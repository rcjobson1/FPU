
module fpu ( clk, rmode, fpu_op, opa, opb, out, inf, snan, qnan, ine, overflow, 
        underflow, zero, div_by_zero );
  input [1:0] rmode;
  input [2:0] fpu_op;
  input [63:0] opa;
  input [63:0] opb;
  output [63:0] out;
  input clk;
  output inf, snan, qnan, ine, overflow, underflow, zero, div_by_zero;
  wire   inf_d, ind_d, qnan_d, snan_d, opa_nan, opb_nan, opa_00, opb_00,
         opa_inf, opb_inf, opb_dn, sign_fasu, nan_sign_d, result_zero_sign_d,
         fasu_op, sign_fasu_r, sign_mul, sign_exe, inf_mul, sign_mul_r,
         inf_mul_r, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265,
         N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276,
         N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287,
         N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298,
         N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, N327,
         N328, N329, N330, N331, N332, N333, N334, N335, N336, N337,
         fract_div_105_, N340, N343, N344, N345, N346, N347, N348, N349, N350,
         N351, N352, N353, N354, N355, N356, N357, N358, N359, N360, N361,
         N362, N363, N364, N365, N366, N367, N368, N369, N370, N371, N372,
         N373, N374, N375, N376, N377, N378, N379, N380, N381, N382, N383,
         N384, N385, N386, N387, N388, N389, N390, N391, N392, N393, N394,
         N395, N396, N501, N502, N503, N504, N505, N506, N507, N508, N509,
         N510, N511, N512, N513, N514, N515, N516, N517, N518, N519, N520,
         N521, N522, N523, N524, N525, N526, N527, N528, N529, N530, N531,
         N532, N533, N534, N535, N536, N537, N538, N539, N540, N541, N542,
         N543, N544, N545, N546, N547, N548, N549, N550, N551, N552, N553,
         N554, N555, N556, N557, N710, N711, N712, N713, N714, N715, N716,
         N717, N718, N719, N720, N721, N722, N723, N724, N725, N726, N727,
         N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738,
         N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749,
         N750, N751, N752, N753, N754, N755, N756, N757, N758, N759, N760,
         N761, N762, N763, N764, N765, N766, N767, N768, N769, opas_r1,
         opas_r2, sign, N789, fasu_op_r1, fasu_op_r2, inf_mul2, N793, N794,
         N795, N796, N797, N798, N799, N800, N801, N802, N803, N804, N805,
         N806, N807, N808, N809, N810, N811, N812, N813, N814, N815, N816,
         N817, N818, N819, N820, N821, N822, N823, N824, N825, N826, N827,
         N828, N829, N830, N831, N832, N833, N834, N835, N836, N837, N838,
         N839, N840, N841, N842, N843, N844, N845, N846, N847, N848, N849,
         N850, N851, N852, N853, N854, N855, N875, N889, N899, N902, N904,
         N906, N911, N912, opa_nan_r, N913, N923, u0_N17, u0_N16, u0_fractb_00,
         u0_fracta_00, u0_expb_00, u0_expa_00, u0_N11, u0_N10, u0_N7, u0_N6,
         u0_snan_r_b, u0_N5, u0_qnan_r_b, u0_snan_r_a, u0_N4, u0_qnan_r_a,
         u0_infb_f_r, u0_infa_f_r, u0_expb_ff, u0_expa_ff, u1_N232, u1_N229,
         u1_fracta_eq_fractb, u1_N220, u1_fracta_lt_fractb, u1_N219, u1_N218,
         u1_add_r, u1_signb_r, u1_signa_r, u1_sign_d, u1_fractb_lt_fracta,
         u1_adj_op_out_sft_0_, u1_adj_op_out_sft_1_, u1_adj_op_out_sft_2_,
         u1_adj_op_out_sft_3_, u1_adj_op_out_sft_4_, u1_adj_op_out_sft_5_,
         u1_adj_op_out_sft_6_, u1_adj_op_out_sft_7_, u1_adj_op_out_sft_8_,
         u1_adj_op_out_sft_9_, u1_adj_op_out_sft_10_, u1_adj_op_out_sft_11_,
         u1_adj_op_out_sft_12_, u1_adj_op_out_sft_13_, u1_adj_op_out_sft_14_,
         u1_adj_op_out_sft_15_, u1_adj_op_out_sft_16_, u1_adj_op_out_sft_17_,
         u1_adj_op_out_sft_18_, u1_adj_op_out_sft_19_, u1_adj_op_out_sft_20_,
         u1_adj_op_out_sft_21_, u1_adj_op_out_sft_22_, u1_adj_op_out_sft_23_,
         u1_adj_op_out_sft_24_, u1_adj_op_out_sft_25_, u1_adj_op_out_sft_26_,
         u1_adj_op_out_sft_27_, u1_adj_op_out_sft_28_, u1_adj_op_out_sft_29_,
         u1_adj_op_out_sft_30_, u1_adj_op_out_sft_31_, u1_adj_op_out_sft_32_,
         u1_adj_op_out_sft_33_, u1_adj_op_out_sft_34_, u1_adj_op_out_sft_35_,
         u1_adj_op_out_sft_36_, u1_adj_op_out_sft_37_, u1_adj_op_out_sft_38_,
         u1_adj_op_out_sft_39_, u1_adj_op_out_sft_40_, u1_adj_op_out_sft_41_,
         u1_adj_op_out_sft_42_, u1_adj_op_out_sft_43_, u1_adj_op_out_sft_44_,
         u1_adj_op_out_sft_45_, u1_adj_op_out_sft_46_, u1_adj_op_out_sft_47_,
         u1_adj_op_out_sft_48_, u1_adj_op_out_sft_49_, u1_adj_op_out_sft_50_,
         u1_adj_op_out_sft_51_, u1_adj_op_out_sft_52_, u1_adj_op_out_sft_53_,
         u1_adj_op_out_sft_54_, u1_adj_op_out_sft_55_, u1_exp_lt_27,
         u1_adj_op_0_, u1_adj_op_3_, u1_adj_op_10_, u1_adj_op_11_,
         u1_adj_op_15_, u1_adj_op_16_, u1_adj_op_17_, u1_adj_op_20_,
         u1_adj_op_21_, u1_adj_op_22_, u1_adj_op_27_, u1_adj_op_28_,
         u1_adj_op_32_, u1_adj_op_36_, u1_adj_op_37_, u1_adj_op_38_,
         u1_adj_op_42_, u1_adj_op_44_, u1_adj_op_51_, u1_N62, u1_N61, u1_N60,
         u1_N59, u1_N58, u1_N57, u1_N56, u1_N55, u1_N54, u1_N53, u1_N52,
         u1_N49, u1_exp_diff_0_, u1_exp_diff_1_, u1_exp_diff_2_,
         u1_exp_diff_3_, u1_exp_diff_4_, u1_exp_diff_5_, u1_exp_diff_6_,
         u1_exp_diff_7_, u1_exp_diff_8_, u1_exp_diff_9_, u1_exp_diff_10_,
         u1_N46, u1_exp_large_0_, u1_exp_large_1_, u1_exp_large_2_,
         u1_exp_large_3_, u1_exp_large_4_, u1_exp_large_5_, u1_exp_large_6_,
         u1_exp_large_7_, u1_exp_large_10_, u1_expa_lt_expb, u2_N157, u2_N121,
         u2_sign_d, u2_N114, u2_N113, u2_N111, u2_exp_ovf_d_0_,
         u2_exp_ovf_d_1_, u2_N86, u2_N85, u2_N84, u2_N83, u2_N82, u2_N81,
         u2_N80, u2_N79, u2_N78, u2_N77, u2_N76, u2_N75, u2_N74, u2_N73,
         u2_N72, u2_N71, u2_N70, u2_N69, u2_N68, u2_N67, u2_N66, u2_N64,
         u2_N63, u2_N62, u2_N61, u2_N60, u2_N59, u2_N58, u2_N57, u2_N56,
         u2_N55, u2_N54, u2_exp_tmp4_1_, u2_exp_tmp4_2_, u2_exp_tmp4_3_,
         u2_exp_tmp4_4_, u2_exp_tmp4_10_, u2_exp_tmp3_0_, u2_exp_tmp3_1_,
         u2_exp_tmp3_2_, u2_exp_tmp3_3_, u2_exp_tmp3_4_, u2_exp_tmp3_5_,
         u2_exp_tmp3_6_, u2_exp_tmp3_7_, u2_exp_tmp3_8_, u2_exp_tmp3_9_,
         u2_exp_tmp3_10_, u2_N53, u2_N52, u2_N51, u2_N50, u2_N49, u2_N48,
         u2_N47, u2_N46, u2_N45, u2_N44, u2_N43, u2_N41, u2_N40, u2_N39,
         u2_N38, u2_N37, u2_N36, u2_N35, u2_N34, u2_N33, u2_N32, u2_N31,
         u2_exp_tmp1_1_, u2_exp_tmp1_2_, u2_exp_tmp1_3_, u2_exp_tmp1_4_,
         u2_N29, u2_N28, u2_N27, u2_N26, u2_N25, u2_N24, u2_N23, u2_N22,
         u2_N21, u2_N20, u2_N19, u2_N18, u2_N17, u2_N16, u2_N15, u2_N14,
         u2_N13, u2_N12, u2_N11, u2_N10, u2_N9, u2_N8, u2_N7, u2_N6, u3_N116,
         u3_N115, u3_N114, u3_N113, u3_N112, u3_N111, u3_N110, u3_N109,
         u3_N108, u3_N107, u3_N106, u3_N105, u3_N104, u3_N103, u3_N102,
         u3_N101, u3_N100, u3_N99, u3_N98, u3_N97, u3_N96, u3_N95, u3_N94,
         u3_N93, u3_N92, u3_N91, u3_N90, u3_N89, u3_N88, u3_N87, u3_N86,
         u3_N85, u3_N84, u3_N83, u3_N82, u3_N81, u3_N80, u3_N79, u3_N78,
         u3_N77, u3_N76, u3_N75, u3_N74, u3_N73, u3_N72, u3_N71, u3_N70,
         u3_N69, u3_N68, u3_N67, u3_N66, u3_N65, u3_N64, u3_N63, u3_N62,
         u3_N61, u3_N60, u3_N59, u3_N58, u3_N57, u3_N56, u3_N55, u3_N54,
         u3_N53, u3_N52, u3_N51, u3_N50, u3_N49, u3_N48, u3_N47, u3_N46,
         u3_N45, u3_N44, u3_N43, u3_N42, u3_N41, u3_N40, u3_N39, u3_N38,
         u3_N37, u3_N36, u3_N35, u3_N34, u3_N33, u3_N32, u3_N31, u3_N30,
         u3_N29, u3_N28, u3_N27, u3_N26, u3_N25, u3_N24, u3_N23, u3_N22,
         u3_N21, u3_N20, u3_N19, u3_N18, u3_N17, u3_N16, u3_N15, u3_N14,
         u3_N13, u3_N12, u3_N11, u3_N10, u3_N9, u3_N8, u3_N7, u3_N6, u3_N5,
         u3_N4, u3_N3, u5_N105, u5_N104, u5_N103, u5_N102, u5_N101, u5_N100,
         u5_N99, u5_N98, u5_N97, u5_N96, u5_N95, u5_N94, u5_N93, u5_N92,
         u5_N91, u5_N90, u5_N89, u5_N88, u5_N87, u5_N86, u5_N85, u5_N84,
         u5_N83, u5_N82, u5_N81, u5_N80, u5_N79, u5_N78, u5_N77, u5_N76,
         u5_N75, u5_N74, u5_N73, u5_N72, u5_N71, u5_N70, u5_N69, u5_N68,
         u5_N67, u5_N66, u5_N65, u5_N64, u5_N63, u5_N62, u5_N61, u5_N60,
         u5_N59, u5_N58, u5_N57, u5_N56, u5_N55, u5_N54, u5_N53, u5_N52,
         u5_N51, u5_N50, u5_N49, u5_N48, u5_N47, u5_N46, u5_N45, u5_N44,
         u5_N43, u5_N42, u5_N41, u5_N40, u5_N39, u5_N38, u5_N37, u5_N36,
         u5_N35, u5_N34, u5_N33, u5_N32, u5_N31, u5_N30, u5_N29, u5_N28,
         u5_N27, u5_N26, u5_N25, u5_N24, u5_N23, u5_N22, u5_N21, u5_N20,
         u5_N19, u5_N18, u5_N17, u5_N16, u5_N15, u5_N14, u5_N13, u5_N12,
         u5_N11, u5_N10, u5_N9, u5_N8, u5_N7, u5_N6, u5_N5, u5_N4, u5_N3,
         u5_N2, u5_N1, u5_N0, u6_N107, u6_N106, u6_N105, u6_N104, u6_N103,
         u6_N102, u6_N101, u6_N100, u6_N99, u6_N98, u6_N97, u6_N96, u6_N95,
         u6_N94, u6_N93, u6_N92, u6_N91, u6_N90, u6_N89, u6_N88, u6_N87,
         u6_N86, u6_N85, u6_N84, u6_N83, u6_N82, u6_N81, u6_N80, u6_N79,
         u6_N78, u6_N77, u6_N76, u6_N75, u6_N74, u6_N73, u6_N72, u6_N71,
         u6_N70, u6_N69, u6_N68, u6_N67, u6_N66, u6_N65, u6_N64, u6_N63,
         u6_N62, u6_N61, u6_N60, u6_N59, u6_N58, u6_N57, u6_N56, u6_N55,
         u6_N52, u6_N51, u6_N50, u6_N49, u6_N48, u6_N47, u6_N46, u6_N45,
         u6_N44, u6_N43, u6_N42, u6_N41, u6_N40, u6_N39, u6_N38, u6_N37,
         u6_N36, u6_N35, u6_N34, u6_N33, u6_N32, u6_N31, u6_N30, u6_N29,
         u6_N28, u6_N27, u6_N26, u6_N25, u6_N24, u6_N23, u6_N22, u6_N21,
         u6_N20, u6_N19, u6_N18, u6_N17, u6_N16, u6_N15, u6_N14, u6_N13,
         u6_N12, u6_N11, u6_N10, u6_N9, u6_N8, u6_N7, u6_N6, u6_N5, u6_N4,
         u6_N3, u6_N2, u6_N1, u6_N0, u4_N6917, u4_N6916, u4_N6915, u4_N6463,
         u4_N6462, u4_N6461, u4_N6460, u4_N6459, u4_N6458, u4_N6457, u4_N6456,
         u4_N6455, u4_N6454, u4_N6410, u4_N6286, u4_N6284, u4_N6283, u4_N6280,
         u4_N6279, u4_N6278, u4_N6251, u4_N6249, u4_N6203, u4_N6194, u4_N6172,
         u4_N6171, u4_div_exp2_0_, u4_div_exp2_1_, u4_div_exp2_2_,
         u4_div_exp2_3_, u4_div_exp2_4_, u4_div_exp2_5_, u4_div_exp2_6_,
         u4_div_exp2_7_, u4_div_exp2_8_, u4_div_exp2_9_, u4_div_exp2_10_,
         u4_div_exp1_0_, u4_div_exp1_1_, u4_div_exp1_2_, u4_div_exp1_3_,
         u4_div_exp1_4_, u4_div_exp1_5_, u4_div_exp1_6_, u4_div_exp1_7_,
         u4_div_exp1_8_, u4_div_exp1_9_, u4_div_exp1_10_, u4_fi_ldz_2a_0_,
         u4_fi_ldz_2a_1_, u4_fi_ldz_2a_2_, u4_fi_ldz_2a_3_, u4_fi_ldz_2a_4_,
         u4_fi_ldz_2a_5_, u4_fi_ldz_2a_6_, u4_ldz_all_0_, u4_ldz_all_1_,
         u4_ldz_all_2_, u4_ldz_all_3_, u4_ldz_all_4_, u4_ldz_all_5_,
         u4_ldz_all_6_, u4_N6142, u4_N6141, u4_N6140, u4_N6139, u4_N6138,
         u4_N6137, u4_N6136, u4_exp_out1_0_, u4_exp_out1_1_, u4_exp_out_pl1_0_,
         u4_exp_out_pl1_1_, u4_exp_out_pl1_2_, u4_exp_out_pl1_3_,
         u4_exp_out_pl1_4_, u4_exp_out_pl1_5_, u4_exp_out_pl1_6_,
         u4_exp_out_pl1_7_, u4_exp_out_pl1_8_, u4_exp_out_pl1_9_,
         u4_exp_out_pl1_10_, u4_fi_ldz_mi1_0_, u4_fi_ldz_mi1_1_,
         u4_fi_ldz_mi1_2_, u4_fi_ldz_mi1_3_, u4_fi_ldz_mi1_4_,
         u4_fi_ldz_mi1_5_, u4_fi_ldz_mi1_6_, u4_N6119, u4_N6118, u4_N6117,
         u4_N6116, u4_N6115, u4_N6114, u4_N6113, u4_N6112, u4_N6111, u4_N6110,
         u4_N6109, u4_N6108, u4_N6107, u4_N6106, u4_N6105, u4_N6104, u4_N6103,
         u4_N6102, u4_N6101, u4_N6100, u4_N6099, u4_N6098, u4_N6097, u4_N6096,
         u4_N6095, u4_N6094, u4_N6093, u4_N6092, u4_N6091, u4_N6090, u4_N6089,
         u4_N6088, u4_N6087, u4_N6086, u4_N6085, u4_N6084, u4_N6083, u4_N6082,
         u4_N6081, u4_N6080, u4_N6079, u4_N6078, u4_N6077, u4_N6076, u4_N6075,
         u4_N6074, u4_N6073, u4_N6072, u4_N6071, u4_N6070, u4_N6069, u4_N6068,
         u4_N6067, u4_N6066, u4_N6065, u4_N6064, u4_N6063, u4_N6062, u4_N6061,
         u4_N6060, u4_N6059, u4_N6058, u4_N6057, u4_N6056, u4_N6055, u4_N6054,
         u4_N6053, u4_N6052, u4_N6051, u4_N6050, u4_N6049, u4_N6048, u4_N6047,
         u4_N6046, u4_N6045, u4_N6044, u4_N6043, u4_N6042, u4_N6041, u4_N6040,
         u4_N6039, u4_N6038, u4_N6037, u4_N6036, u4_N6035, u4_N6034, u4_N6033,
         u4_N6032, u4_N6031, u4_N6030, u4_N6029, u4_N6028, u4_N6027, u4_N6026,
         u4_N6025, u4_N6024, u4_N6023, u4_N6022, u4_N6021, u4_N6020, u4_N6019,
         u4_N6018, u4_N6017, u4_N6016, u4_N6015, u4_N6014, u4_N6011, u4_N6010,
         u4_N6009, u4_N6008, u4_N6007, u4_N6006, u4_N6005, u4_N6004, u4_N6003,
         u4_N6002, u4_N6001, u4_N6000, u4_N5999, u4_N5998, u4_N5997, u4_N5996,
         u4_N5995, u4_N5994, u4_N5993, u4_N5992, u4_N5991, u4_N5990, u4_N5989,
         u4_N5988, u4_N5987, u4_N5986, u4_N5985, u4_N5984, u4_N5983, u4_N5982,
         u4_N5981, u4_N5980, u4_N5979, u4_N5978, u4_N5977, u4_N5976, u4_N5975,
         u4_N5974, u4_N5973, u4_N5972, u4_N5971, u4_N5970, u4_N5969, u4_N5968,
         u4_N5967, u4_N5966, u4_N5965, u4_N5964, u4_N5963, u4_N5962, u4_N5961,
         u4_N5960, u4_N5959, u4_N5958, u4_N5957, u4_N5956, u4_N5955, u4_N5954,
         u4_N5953, u4_N5952, u4_N5951, u4_N5950, u4_N5949, u4_N5948, u4_N5947,
         u4_N5946, u4_N5945, u4_N5944, u4_N5943, u4_N5942, u4_N5941, u4_N5940,
         u4_N5939, u4_N5938, u4_N5937, u4_N5936, u4_N5935, u4_N5934, u4_N5933,
         u4_N5932, u4_N5931, u4_N5930, u4_N5929, u4_N5928, u4_N5927, u4_N5926,
         u4_N5925, u4_N5924, u4_N5923, u4_N5922, u4_N5921, u4_N5920, u4_N5919,
         u4_N5918, u4_N5917, u4_N5916, u4_N5915, u4_N5914, u4_N5913, u4_N5912,
         u4_N5911, u4_N5910, u4_N5909, u4_N5908, u4_N5907, u4_N5906, u4_N5904,
         u4_exp_in_pl1_0_, u4_exp_in_pl1_1_, u4_exp_in_pl1_2_,
         u4_exp_in_pl1_3_, u4_exp_in_pl1_4_, u4_exp_in_pl1_5_,
         u4_exp_in_pl1_6_, u4_exp_in_pl1_7_, u4_exp_in_pl1_8_,
         u4_exp_in_pl1_9_, u4_exp_in_pl1_10_, u4_exp_in_pl1_11_,
         u4_f2i_shft_1_, u4_f2i_shft_2_, u4_f2i_shft_3_, u4_f2i_shft_4_,
         u4_f2i_shft_5_, u4_f2i_shft_6_, u4_f2i_shft_7_, u4_f2i_shft_8_,
         u4_f2i_shft_9_, u4_f2i_shft_10_, u4_N5843, u4_div_shft3_0_,
         u4_div_shft3_1_, u4_div_shft3_2_, u4_div_shft3_3_, u4_div_shft3_4_,
         u4_div_shft3_5_, u4_div_shft3_6_, u4_div_shft3_7_, u4_div_shft3_8_,
         u4_div_shft3_9_, u4_div_shft3_10_, u4_exp_in_mi1_1_, u4_exp_in_mi1_2_,
         u4_exp_in_mi1_3_, u4_exp_in_mi1_4_, u4_exp_in_mi1_5_,
         u4_exp_in_mi1_6_, u4_exp_in_mi1_7_, u4_exp_in_mi1_8_,
         u4_exp_in_mi1_9_, u4_exp_in_mi1_10_, u4_exp_in_mi1_11_, u4_N5837,
         u4_N5836, u4_fract_out_pl1_0_, u4_fract_out_pl1_1_,
         u4_fract_out_pl1_2_, u4_fract_out_pl1_3_, u4_fract_out_pl1_4_,
         u4_fract_out_pl1_5_, u4_fract_out_pl1_6_, u4_fract_out_pl1_7_,
         u4_fract_out_pl1_8_, u4_fract_out_pl1_9_, u4_fract_out_pl1_10_,
         u4_fract_out_pl1_11_, u4_fract_out_pl1_12_, u4_fract_out_pl1_13_,
         u4_fract_out_pl1_14_, u4_fract_out_pl1_15_, u4_fract_out_pl1_16_,
         u4_fract_out_pl1_17_, u4_fract_out_pl1_18_, u4_fract_out_pl1_19_,
         u4_fract_out_pl1_20_, u4_fract_out_pl1_21_, u4_fract_out_pl1_22_,
         u4_fract_out_pl1_23_, u4_fract_out_pl1_24_, u4_fract_out_pl1_25_,
         u4_fract_out_pl1_26_, u4_fract_out_pl1_27_, u4_fract_out_pl1_28_,
         u4_fract_out_pl1_29_, u4_fract_out_pl1_30_, u4_fract_out_pl1_31_,
         u4_fract_out_pl1_32_, u4_fract_out_pl1_33_, u4_fract_out_pl1_34_,
         u4_fract_out_pl1_35_, u4_fract_out_pl1_36_, u4_fract_out_pl1_37_,
         u4_fract_out_pl1_38_, u4_fract_out_pl1_39_, u4_fract_out_pl1_40_,
         u4_fract_out_pl1_41_, u4_fract_out_pl1_42_, u4_fract_out_pl1_43_,
         u4_fract_out_pl1_44_, u4_fract_out_pl1_45_, u4_fract_out_pl1_46_,
         u4_fract_out_pl1_47_, u4_fract_out_pl1_48_, u4_fract_out_pl1_49_,
         u4_fract_out_pl1_50_, u4_fract_out_pl1_51_, u4_fract_out_pl1_52_,
         u4_exp_next_mi_0_, u4_exp_next_mi_1_, u4_exp_next_mi_2_,
         u4_exp_next_mi_3_, u4_exp_next_mi_4_, u4_exp_next_mi_5_,
         u4_exp_next_mi_6_, u4_exp_next_mi_7_, u4_exp_next_mi_8_,
         u4_exp_next_mi_9_, u4_exp_next_mi_10_, u4_exp_next_mi_11_,
         u4_fract_out_0_, u4_fract_out_1_, u4_fract_out_2_, u4_fract_out_3_,
         u4_fract_out_4_, u4_fract_out_5_, u4_fract_out_6_, u4_fract_out_7_,
         u4_fract_out_8_, u4_fract_out_9_, u4_fract_out_10_, u4_fract_out_11_,
         u4_fract_out_12_, u4_fract_out_13_, u4_fract_out_14_,
         u4_fract_out_15_, u4_fract_out_16_, u4_fract_out_17_,
         u4_fract_out_18_, u4_fract_out_19_, u4_fract_out_20_,
         u4_fract_out_21_, u4_fract_out_22_, u4_fract_out_23_,
         u4_fract_out_24_, u4_fract_out_25_, u4_fract_out_26_,
         u4_fract_out_27_, u4_fract_out_28_, u4_fract_out_29_,
         u4_fract_out_30_, u4_fract_out_31_, u4_fract_out_32_,
         u4_fract_out_33_, u4_fract_out_34_, u4_fract_out_35_,
         u4_fract_out_36_, u4_fract_out_37_, u4_fract_out_38_,
         u4_fract_out_39_, u4_fract_out_40_, u4_fract_out_41_,
         u4_fract_out_42_, u4_fract_out_43_, u4_fract_out_44_,
         u4_fract_out_45_, u4_fract_out_46_, u4_fract_out_47_,
         u4_fract_out_48_, u4_fract_out_49_, u4_fract_out_50_,
         u4_fract_out_51_, u4_exp_out_0_, u4_exp_out_1_, u4_exp_out_2_,
         u4_exp_out_3_, u4_exp_out_4_, u4_exp_out_5_, u4_exp_out_6_,
         u4_exp_out_7_, u4_exp_out_8_, u4_exp_out_9_, u4_exp_out_10_,
         u4_fi_ldz_1_, u4_fi_ldz_2_, u4_fi_ldz_3_, u4_fi_ldz_4_, u4_fi_ldz_5_,
         u4_fi_ldz_6_, n203, n204, n205, n2388, n2389, n2390, n2391, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3621, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4194, n4195, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, u4_ldz_dif_9_, u4_ldz_dif_8_,
         u4_ldz_dif_7_, u4_ldz_dif_6_, u4_ldz_dif_5_, u4_ldz_dif_4_,
         u4_ldz_dif_3_, u4_ldz_dif_2_, u4_ldz_dif_1_, u4_ldz_dif_10_,
         u4_ldz_dif_0_, u2_lt_135_A_0_, u2_lt_135_A_5_, u2_lt_135_A_6_,
         u2_lt_135_A_7_, u2_lt_135_A_8_, u2_lt_135_A_9_, u2_gt_145_B_11_,
         u4_sub_463_carry_2_, u4_sub_463_carry_3_, u4_sub_463_carry_4_,
         u4_sub_463_carry_5_, u4_sub_463_carry_6_, u4_sub_468_A_2_,
         u4_sub_468_A_3_, u4_sub_468_A_4_, u4_sub_468_A_5_, u4_sub_468_A_7_,
         u4_sub_468_A_9_, u4_sub_468_A_10_, u4_sub_417_carry_2_,
         u4_sub_417_carry_3_, u4_sub_417_carry_4_, u4_sub_417_carry_5_,
         u4_sub_417_carry_6_, u4_sub_417_carry_7_, u4_sub_417_carry_8_,
         u4_sub_417_carry_9_, u4_sub_417_carry_10_, u2_sub_116_carry_2_,
         u2_sub_116_carry_3_, u2_sub_116_carry_4_, u2_sub_116_carry_5_,
         u2_sub_116_carry_6_, u2_sub_116_carry_7_, u2_sub_116_carry_8_,
         u2_sub_116_carry_9_, u2_sub_116_carry_10_, u2_sub_116_carry_11_,
         u2_add_116_carry_2_, u2_add_116_carry_3_, u2_add_116_carry_4_,
         u2_add_116_carry_5_, u2_add_116_carry_6_, u2_add_116_carry_7_,
         u2_add_116_carry_8_, u2_add_116_carry_9_, u2_add_116_carry_10_,
         u2_add_116_carry_11_, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, u4_sub_473_n14, u4_sub_473_n13, u4_sub_473_n12,
         u4_sub_473_n11, u4_sub_473_n10, u4_sub_473_n9, u4_sub_473_n8,
         u4_sub_473_n7, u4_sub_473_n6, u4_sub_473_n5, u4_sub_473_n4,
         u4_sub_473_n3, u4_sub_473_n2, u4_sub_473_n1, u4_sub_473_carry_1_,
         u4_sub_473_carry_2_, u4_sub_473_carry_3_, u4_sub_473_carry_4_,
         u4_sub_473_carry_5_, u4_sub_473_carry_6_, u4_sub_473_carry_7_,
         u4_sub_473_carry_8_, u4_sub_473_carry_9_, u4_sub_473_carry_10_,
         u4_sub_472_n14, u4_sub_472_n13, u4_sub_472_n12, u4_sub_472_n11,
         u4_sub_472_n10, u4_sub_472_n9, u4_sub_472_n8, u4_sub_472_n7,
         u4_sub_472_n6, u4_sub_472_n5, u4_sub_472_n4, u4_sub_472_n3,
         u4_sub_472_n2, u4_sub_472_n1, u4_sub_472_carry_1_,
         u4_sub_472_carry_2_, u4_sub_472_carry_3_, u4_sub_472_carry_4_,
         u4_sub_472_carry_5_, u4_sub_472_carry_6_, u4_sub_472_carry_7_,
         u4_sub_472_carry_8_, u4_sub_472_carry_9_, u4_sub_472_carry_10_,
         u4_sll_454_n88, u4_sll_454_n87, u4_sll_454_n86, u4_sll_454_n85,
         u4_sll_454_n84, u4_sll_454_n83, u4_sll_454_n82, u4_sll_454_n81,
         u4_sll_454_n80, u4_sll_454_n79, u4_sll_454_n78, u4_sll_454_n77,
         u4_sll_454_n76, u4_sll_454_n75, u4_sll_454_n74, u4_sll_454_n73,
         u4_sll_454_n72, u4_sll_454_n71, u4_sll_454_n70, u4_sll_454_n69,
         u4_sll_454_n68, u4_sll_454_n67, u4_sll_454_n66, u4_sll_454_n65,
         u4_sll_454_n64, u4_sll_454_n63, u4_sll_454_n62, u4_sll_454_n61,
         u4_sll_454_n60, u4_sll_454_n59, u4_sll_454_n58, u4_sll_454_n57,
         u4_sll_454_n56, u4_sll_454_n55, u4_sll_454_n54, u4_sll_454_n53,
         u4_sll_454_n52, u4_sll_454_n51, u4_sll_454_n50, u4_sll_454_n49,
         u4_sll_454_n48, u4_sll_454_n47, u4_sll_454_n46, u4_sll_454_n45,
         u4_sll_454_n44, u4_sll_454_n43, u4_sll_454_n42, u4_sll_454_n41,
         u4_sll_454_n40, u4_sll_454_n39, u4_sll_454_n38, u4_sll_454_n37,
         u4_sll_454_n36, u4_sll_454_n35, u4_sll_454_n34, u4_sll_454_n33,
         u4_sll_454_n32, u4_sll_454_n31, u4_sll_454_n30, u4_sll_454_n29,
         u4_sll_454_n28, u4_sll_454_n27, u4_sll_454_n26, u4_sll_454_n25,
         u4_sll_454_n24, u4_sll_454_n23, u4_sll_454_n22, u4_sll_454_n21,
         u4_sll_454_n20, u4_sll_454_n19, u4_sll_454_n18, u4_sll_454_n17,
         u4_sll_454_n16, u4_sll_454_n15, u4_sll_454_n14, u4_sll_454_n13,
         u4_sll_454_n12, u4_sll_454_n11, u4_sll_454_n10, u4_sll_454_n9,
         u4_sll_454_n8, u4_sll_454_n7, u4_sll_454_n6, u4_sll_454_n5,
         u4_sll_454_n4, u4_sll_454_n3, u4_sll_454_n2, u4_sll_454_n1,
         u4_sll_454_ML_int_7__64_, u4_sll_454_ML_int_7__65_,
         u4_sll_454_ML_int_7__66_, u4_sll_454_ML_int_7__67_,
         u4_sll_454_ML_int_7__68_, u4_sll_454_ML_int_7__69_,
         u4_sll_454_ML_int_7__70_, u4_sll_454_ML_int_7__71_,
         u4_sll_454_ML_int_7__72_, u4_sll_454_ML_int_7__73_,
         u4_sll_454_ML_int_7__74_, u4_sll_454_ML_int_7__75_,
         u4_sll_454_ML_int_7__76_, u4_sll_454_ML_int_7__77_,
         u4_sll_454_ML_int_7__78_, u4_sll_454_ML_int_7__79_,
         u4_sll_454_ML_int_7__80_, u4_sll_454_ML_int_7__81_,
         u4_sll_454_ML_int_7__82_, u4_sll_454_ML_int_7__83_,
         u4_sll_454_ML_int_7__84_, u4_sll_454_ML_int_7__85_,
         u4_sll_454_ML_int_7__86_, u4_sll_454_ML_int_7__87_,
         u4_sll_454_ML_int_7__88_, u4_sll_454_ML_int_7__89_,
         u4_sll_454_ML_int_7__90_, u4_sll_454_ML_int_7__91_,
         u4_sll_454_ML_int_7__92_, u4_sll_454_ML_int_7__93_,
         u4_sll_454_ML_int_7__94_, u4_sll_454_ML_int_7__95_,
         u4_sll_454_ML_int_7__96_, u4_sll_454_ML_int_7__97_,
         u4_sll_454_ML_int_7__98_, u4_sll_454_ML_int_7__99_,
         u4_sll_454_ML_int_7__100_, u4_sll_454_ML_int_7__101_,
         u4_sll_454_ML_int_7__102_, u4_sll_454_ML_int_7__103_,
         u4_sll_454_ML_int_7__104_, u4_sll_454_ML_int_7__105_,
         u4_sll_454_ML_int_6__0_, u4_sll_454_ML_int_6__1_,
         u4_sll_454_ML_int_6__2_, u4_sll_454_ML_int_6__3_,
         u4_sll_454_ML_int_6__4_, u4_sll_454_ML_int_6__5_,
         u4_sll_454_ML_int_6__6_, u4_sll_454_ML_int_6__7_,
         u4_sll_454_ML_int_6__8_, u4_sll_454_ML_int_6__9_,
         u4_sll_454_ML_int_6__10_, u4_sll_454_ML_int_6__11_,
         u4_sll_454_ML_int_6__12_, u4_sll_454_ML_int_6__13_,
         u4_sll_454_ML_int_6__14_, u4_sll_454_ML_int_6__15_,
         u4_sll_454_ML_int_6__16_, u4_sll_454_ML_int_6__17_,
         u4_sll_454_ML_int_6__18_, u4_sll_454_ML_int_6__19_,
         u4_sll_454_ML_int_6__20_, u4_sll_454_ML_int_6__21_,
         u4_sll_454_ML_int_6__22_, u4_sll_454_ML_int_6__23_,
         u4_sll_454_ML_int_6__24_, u4_sll_454_ML_int_6__25_,
         u4_sll_454_ML_int_6__26_, u4_sll_454_ML_int_6__27_,
         u4_sll_454_ML_int_6__28_, u4_sll_454_ML_int_6__29_,
         u4_sll_454_ML_int_6__30_, u4_sll_454_ML_int_6__31_,
         u4_sll_454_ML_int_6__32_, u4_sll_454_ML_int_6__33_,
         u4_sll_454_ML_int_6__34_, u4_sll_454_ML_int_6__35_,
         u4_sll_454_ML_int_6__36_, u4_sll_454_ML_int_6__37_,
         u4_sll_454_ML_int_6__38_, u4_sll_454_ML_int_6__39_,
         u4_sll_454_ML_int_6__40_, u4_sll_454_ML_int_6__41_,
         u4_sll_454_ML_int_6__42_, u4_sll_454_ML_int_6__43_,
         u4_sll_454_ML_int_6__44_, u4_sll_454_ML_int_6__45_,
         u4_sll_454_ML_int_6__46_, u4_sll_454_ML_int_6__47_,
         u4_sll_454_ML_int_6__48_, u4_sll_454_ML_int_6__49_,
         u4_sll_454_ML_int_6__50_, u4_sll_454_ML_int_6__51_,
         u4_sll_454_ML_int_6__52_, u4_sll_454_ML_int_6__53_,
         u4_sll_454_ML_int_6__54_, u4_sll_454_ML_int_6__55_,
         u4_sll_454_ML_int_6__56_, u4_sll_454_ML_int_6__57_,
         u4_sll_454_ML_int_6__58_, u4_sll_454_ML_int_6__59_,
         u4_sll_454_ML_int_6__60_, u4_sll_454_ML_int_6__61_,
         u4_sll_454_ML_int_6__62_, u4_sll_454_ML_int_6__63_,
         u4_sll_454_ML_int_6__64_, u4_sll_454_ML_int_6__65_,
         u4_sll_454_ML_int_6__66_, u4_sll_454_ML_int_6__67_,
         u4_sll_454_ML_int_6__68_, u4_sll_454_ML_int_6__69_,
         u4_sll_454_ML_int_6__70_, u4_sll_454_ML_int_6__71_,
         u4_sll_454_ML_int_6__72_, u4_sll_454_ML_int_6__73_,
         u4_sll_454_ML_int_6__74_, u4_sll_454_ML_int_6__75_,
         u4_sll_454_ML_int_6__76_, u4_sll_454_ML_int_6__77_,
         u4_sll_454_ML_int_6__78_, u4_sll_454_ML_int_6__79_,
         u4_sll_454_ML_int_6__80_, u4_sll_454_ML_int_6__81_,
         u4_sll_454_ML_int_6__82_, u4_sll_454_ML_int_6__83_,
         u4_sll_454_ML_int_6__84_, u4_sll_454_ML_int_6__85_,
         u4_sll_454_ML_int_6__86_, u4_sll_454_ML_int_6__87_,
         u4_sll_454_ML_int_6__88_, u4_sll_454_ML_int_6__89_,
         u4_sll_454_ML_int_6__90_, u4_sll_454_ML_int_6__91_,
         u4_sll_454_ML_int_6__92_, u4_sll_454_ML_int_6__93_,
         u4_sll_454_ML_int_6__94_, u4_sll_454_ML_int_6__95_,
         u4_sll_454_ML_int_6__96_, u4_sll_454_ML_int_6__97_,
         u4_sll_454_ML_int_6__98_, u4_sll_454_ML_int_6__99_,
         u4_sll_454_ML_int_6__100_, u4_sll_454_ML_int_6__101_,
         u4_sll_454_ML_int_6__102_, u4_sll_454_ML_int_6__103_,
         u4_sll_454_ML_int_6__104_, u4_sll_454_ML_int_6__105_,
         u4_sll_454_ML_int_5__0_, u4_sll_454_ML_int_5__1_,
         u4_sll_454_ML_int_5__2_, u4_sll_454_ML_int_5__3_,
         u4_sll_454_ML_int_5__4_, u4_sll_454_ML_int_5__5_,
         u4_sll_454_ML_int_5__6_, u4_sll_454_ML_int_5__7_,
         u4_sll_454_ML_int_5__8_, u4_sll_454_ML_int_5__9_,
         u4_sll_454_ML_int_5__10_, u4_sll_454_ML_int_5__11_,
         u4_sll_454_ML_int_5__12_, u4_sll_454_ML_int_5__13_,
         u4_sll_454_ML_int_5__14_, u4_sll_454_ML_int_5__15_,
         u4_sll_454_ML_int_5__16_, u4_sll_454_ML_int_5__17_,
         u4_sll_454_ML_int_5__18_, u4_sll_454_ML_int_5__19_,
         u4_sll_454_ML_int_5__20_, u4_sll_454_ML_int_5__21_,
         u4_sll_454_ML_int_5__22_, u4_sll_454_ML_int_5__23_,
         u4_sll_454_ML_int_5__24_, u4_sll_454_ML_int_5__25_,
         u4_sll_454_ML_int_5__26_, u4_sll_454_ML_int_5__27_,
         u4_sll_454_ML_int_5__28_, u4_sll_454_ML_int_5__29_,
         u4_sll_454_ML_int_5__30_, u4_sll_454_ML_int_5__31_,
         u4_sll_454_ML_int_5__32_, u4_sll_454_ML_int_5__33_,
         u4_sll_454_ML_int_5__34_, u4_sll_454_ML_int_5__35_,
         u4_sll_454_ML_int_5__36_, u4_sll_454_ML_int_5__37_,
         u4_sll_454_ML_int_5__38_, u4_sll_454_ML_int_5__39_,
         u4_sll_454_ML_int_5__40_, u4_sll_454_ML_int_5__41_,
         u4_sll_454_ML_int_5__42_, u4_sll_454_ML_int_5__43_,
         u4_sll_454_ML_int_5__44_, u4_sll_454_ML_int_5__45_,
         u4_sll_454_ML_int_5__46_, u4_sll_454_ML_int_5__47_,
         u4_sll_454_ML_int_5__48_, u4_sll_454_ML_int_5__49_,
         u4_sll_454_ML_int_5__50_, u4_sll_454_ML_int_5__51_,
         u4_sll_454_ML_int_5__52_, u4_sll_454_ML_int_5__53_,
         u4_sll_454_ML_int_5__54_, u4_sll_454_ML_int_5__55_,
         u4_sll_454_ML_int_5__56_, u4_sll_454_ML_int_5__57_,
         u4_sll_454_ML_int_5__58_, u4_sll_454_ML_int_5__59_,
         u4_sll_454_ML_int_5__60_, u4_sll_454_ML_int_5__61_,
         u4_sll_454_ML_int_5__62_, u4_sll_454_ML_int_5__63_,
         u4_sll_454_ML_int_5__64_, u4_sll_454_ML_int_5__65_,
         u4_sll_454_ML_int_5__66_, u4_sll_454_ML_int_5__67_,
         u4_sll_454_ML_int_5__68_, u4_sll_454_ML_int_5__69_,
         u4_sll_454_ML_int_5__70_, u4_sll_454_ML_int_5__71_,
         u4_sll_454_ML_int_5__72_, u4_sll_454_ML_int_5__73_,
         u4_sll_454_ML_int_5__74_, u4_sll_454_ML_int_5__75_,
         u4_sll_454_ML_int_5__76_, u4_sll_454_ML_int_5__77_,
         u4_sll_454_ML_int_5__78_, u4_sll_454_ML_int_5__79_,
         u4_sll_454_ML_int_5__80_, u4_sll_454_ML_int_5__81_,
         u4_sll_454_ML_int_5__82_, u4_sll_454_ML_int_5__83_,
         u4_sll_454_ML_int_5__84_, u4_sll_454_ML_int_5__85_,
         u4_sll_454_ML_int_5__86_, u4_sll_454_ML_int_5__87_,
         u4_sll_454_ML_int_5__88_, u4_sll_454_ML_int_5__89_,
         u4_sll_454_ML_int_5__90_, u4_sll_454_ML_int_5__91_,
         u4_sll_454_ML_int_5__92_, u4_sll_454_ML_int_5__93_,
         u4_sll_454_ML_int_5__94_, u4_sll_454_ML_int_5__95_,
         u4_sll_454_ML_int_5__96_, u4_sll_454_ML_int_5__97_,
         u4_sll_454_ML_int_5__98_, u4_sll_454_ML_int_5__99_,
         u4_sll_454_ML_int_5__100_, u4_sll_454_ML_int_5__101_,
         u4_sll_454_ML_int_5__102_, u4_sll_454_ML_int_5__103_,
         u4_sll_454_ML_int_5__104_, u4_sll_454_ML_int_5__105_,
         u4_sll_454_ML_int_4__0_, u4_sll_454_ML_int_4__1_,
         u4_sll_454_ML_int_4__2_, u4_sll_454_ML_int_4__3_,
         u4_sll_454_ML_int_4__4_, u4_sll_454_ML_int_4__5_,
         u4_sll_454_ML_int_4__6_, u4_sll_454_ML_int_4__7_,
         u4_sll_454_ML_int_4__8_, u4_sll_454_ML_int_4__9_,
         u4_sll_454_ML_int_4__10_, u4_sll_454_ML_int_4__11_,
         u4_sll_454_ML_int_4__12_, u4_sll_454_ML_int_4__13_,
         u4_sll_454_ML_int_4__14_, u4_sll_454_ML_int_4__15_,
         u4_sll_454_ML_int_4__16_, u4_sll_454_ML_int_4__17_,
         u4_sll_454_ML_int_4__18_, u4_sll_454_ML_int_4__19_,
         u4_sll_454_ML_int_4__20_, u4_sll_454_ML_int_4__21_,
         u4_sll_454_ML_int_4__22_, u4_sll_454_ML_int_4__23_,
         u4_sll_454_ML_int_4__24_, u4_sll_454_ML_int_4__25_,
         u4_sll_454_ML_int_4__26_, u4_sll_454_ML_int_4__27_,
         u4_sll_454_ML_int_4__28_, u4_sll_454_ML_int_4__29_,
         u4_sll_454_ML_int_4__30_, u4_sll_454_ML_int_4__31_,
         u4_sll_454_ML_int_4__32_, u4_sll_454_ML_int_4__33_,
         u4_sll_454_ML_int_4__34_, u4_sll_454_ML_int_4__35_,
         u4_sll_454_ML_int_4__36_, u4_sll_454_ML_int_4__37_,
         u4_sll_454_ML_int_4__38_, u4_sll_454_ML_int_4__39_,
         u4_sll_454_ML_int_4__40_, u4_sll_454_ML_int_4__41_,
         u4_sll_454_ML_int_4__42_, u4_sll_454_ML_int_4__43_,
         u4_sll_454_ML_int_4__44_, u4_sll_454_ML_int_4__45_,
         u4_sll_454_ML_int_4__46_, u4_sll_454_ML_int_4__47_,
         u4_sll_454_ML_int_4__48_, u4_sll_454_ML_int_4__49_,
         u4_sll_454_ML_int_4__50_, u4_sll_454_ML_int_4__51_,
         u4_sll_454_ML_int_4__52_, u4_sll_454_ML_int_4__53_,
         u4_sll_454_ML_int_4__54_, u4_sll_454_ML_int_4__55_,
         u4_sll_454_ML_int_4__56_, u4_sll_454_ML_int_4__57_,
         u4_sll_454_ML_int_4__58_, u4_sll_454_ML_int_4__59_,
         u4_sll_454_ML_int_4__60_, u4_sll_454_ML_int_4__61_,
         u4_sll_454_ML_int_4__62_, u4_sll_454_ML_int_4__63_,
         u4_sll_454_ML_int_4__64_, u4_sll_454_ML_int_4__65_,
         u4_sll_454_ML_int_4__66_, u4_sll_454_ML_int_4__67_,
         u4_sll_454_ML_int_4__68_, u4_sll_454_ML_int_4__69_,
         u4_sll_454_ML_int_4__70_, u4_sll_454_ML_int_4__71_,
         u4_sll_454_ML_int_4__72_, u4_sll_454_ML_int_4__73_,
         u4_sll_454_ML_int_4__74_, u4_sll_454_ML_int_4__75_,
         u4_sll_454_ML_int_4__76_, u4_sll_454_ML_int_4__77_,
         u4_sll_454_ML_int_4__78_, u4_sll_454_ML_int_4__79_,
         u4_sll_454_ML_int_4__80_, u4_sll_454_ML_int_4__81_,
         u4_sll_454_ML_int_4__82_, u4_sll_454_ML_int_4__83_,
         u4_sll_454_ML_int_4__84_, u4_sll_454_ML_int_4__85_,
         u4_sll_454_ML_int_4__86_, u4_sll_454_ML_int_4__87_,
         u4_sll_454_ML_int_4__88_, u4_sll_454_ML_int_4__89_,
         u4_sll_454_ML_int_4__90_, u4_sll_454_ML_int_4__91_,
         u4_sll_454_ML_int_4__92_, u4_sll_454_ML_int_4__93_,
         u4_sll_454_ML_int_4__94_, u4_sll_454_ML_int_4__95_,
         u4_sll_454_ML_int_4__96_, u4_sll_454_ML_int_4__97_,
         u4_sll_454_ML_int_4__98_, u4_sll_454_ML_int_4__99_,
         u4_sll_454_ML_int_4__100_, u4_sll_454_ML_int_4__101_,
         u4_sll_454_ML_int_4__102_, u4_sll_454_ML_int_4__103_,
         u4_sll_454_ML_int_4__104_, u4_sll_454_ML_int_4__105_,
         u4_sll_454_ML_int_3__0_, u4_sll_454_ML_int_3__1_,
         u4_sll_454_ML_int_3__2_, u4_sll_454_ML_int_3__3_,
         u4_sll_454_ML_int_3__4_, u4_sll_454_ML_int_3__5_,
         u4_sll_454_ML_int_3__6_, u4_sll_454_ML_int_3__7_,
         u4_sll_454_ML_int_3__8_, u4_sll_454_ML_int_3__9_,
         u4_sll_454_ML_int_3__10_, u4_sll_454_ML_int_3__11_,
         u4_sll_454_ML_int_3__12_, u4_sll_454_ML_int_3__13_,
         u4_sll_454_ML_int_3__14_, u4_sll_454_ML_int_3__15_,
         u4_sll_454_ML_int_3__16_, u4_sll_454_ML_int_3__17_,
         u4_sll_454_ML_int_3__18_, u4_sll_454_ML_int_3__19_,
         u4_sll_454_ML_int_3__20_, u4_sll_454_ML_int_3__21_,
         u4_sll_454_ML_int_3__22_, u4_sll_454_ML_int_3__23_,
         u4_sll_454_ML_int_3__24_, u4_sll_454_ML_int_3__25_,
         u4_sll_454_ML_int_3__26_, u4_sll_454_ML_int_3__27_,
         u4_sll_454_ML_int_3__28_, u4_sll_454_ML_int_3__29_,
         u4_sll_454_ML_int_3__30_, u4_sll_454_ML_int_3__31_,
         u4_sll_454_ML_int_3__32_, u4_sll_454_ML_int_3__33_,
         u4_sll_454_ML_int_3__34_, u4_sll_454_ML_int_3__35_,
         u4_sll_454_ML_int_3__36_, u4_sll_454_ML_int_3__37_,
         u4_sll_454_ML_int_3__38_, u4_sll_454_ML_int_3__39_,
         u4_sll_454_ML_int_3__40_, u4_sll_454_ML_int_3__41_,
         u4_sll_454_ML_int_3__42_, u4_sll_454_ML_int_3__43_,
         u4_sll_454_ML_int_3__44_, u4_sll_454_ML_int_3__45_,
         u4_sll_454_ML_int_3__46_, u4_sll_454_ML_int_3__47_,
         u4_sll_454_ML_int_3__48_, u4_sll_454_ML_int_3__49_,
         u4_sll_454_ML_int_3__50_, u4_sll_454_ML_int_3__51_,
         u4_sll_454_ML_int_3__52_, u4_sll_454_ML_int_3__53_,
         u4_sll_454_ML_int_3__54_, u4_sll_454_ML_int_3__55_,
         u4_sll_454_ML_int_3__56_, u4_sll_454_ML_int_3__57_,
         u4_sll_454_ML_int_3__58_, u4_sll_454_ML_int_3__59_,
         u4_sll_454_ML_int_3__60_, u4_sll_454_ML_int_3__61_,
         u4_sll_454_ML_int_3__62_, u4_sll_454_ML_int_3__63_,
         u4_sll_454_ML_int_3__64_, u4_sll_454_ML_int_3__65_,
         u4_sll_454_ML_int_3__66_, u4_sll_454_ML_int_3__67_,
         u4_sll_454_ML_int_3__68_, u4_sll_454_ML_int_3__69_,
         u4_sll_454_ML_int_3__70_, u4_sll_454_ML_int_3__71_,
         u4_sll_454_ML_int_3__72_, u4_sll_454_ML_int_3__73_,
         u4_sll_454_ML_int_3__74_, u4_sll_454_ML_int_3__75_,
         u4_sll_454_ML_int_3__76_, u4_sll_454_ML_int_3__77_,
         u4_sll_454_ML_int_3__78_, u4_sll_454_ML_int_3__79_,
         u4_sll_454_ML_int_3__80_, u4_sll_454_ML_int_3__81_,
         u4_sll_454_ML_int_3__82_, u4_sll_454_ML_int_3__83_,
         u4_sll_454_ML_int_3__84_, u4_sll_454_ML_int_3__85_,
         u4_sll_454_ML_int_3__86_, u4_sll_454_ML_int_3__87_,
         u4_sll_454_ML_int_3__88_, u4_sll_454_ML_int_3__89_,
         u4_sll_454_ML_int_3__90_, u4_sll_454_ML_int_3__91_,
         u4_sll_454_ML_int_3__92_, u4_sll_454_ML_int_3__93_,
         u4_sll_454_ML_int_3__94_, u4_sll_454_ML_int_3__95_,
         u4_sll_454_ML_int_3__96_, u4_sll_454_ML_int_3__97_,
         u4_sll_454_ML_int_3__98_, u4_sll_454_ML_int_3__99_,
         u4_sll_454_ML_int_3__100_, u4_sll_454_ML_int_3__101_,
         u4_sll_454_ML_int_3__102_, u4_sll_454_ML_int_3__103_,
         u4_sll_454_ML_int_3__104_, u4_sll_454_ML_int_3__105_,
         u4_sll_454_ML_int_2__0_, u4_sll_454_ML_int_2__1_,
         u4_sll_454_ML_int_2__2_, u4_sll_454_ML_int_2__3_,
         u4_sll_454_ML_int_2__4_, u4_sll_454_ML_int_2__5_,
         u4_sll_454_ML_int_2__6_, u4_sll_454_ML_int_2__7_,
         u4_sll_454_ML_int_2__8_, u4_sll_454_ML_int_2__9_,
         u4_sll_454_ML_int_2__10_, u4_sll_454_ML_int_2__11_,
         u4_sll_454_ML_int_2__12_, u4_sll_454_ML_int_2__13_,
         u4_sll_454_ML_int_2__14_, u4_sll_454_ML_int_2__15_,
         u4_sll_454_ML_int_2__16_, u4_sll_454_ML_int_2__17_,
         u4_sll_454_ML_int_2__18_, u4_sll_454_ML_int_2__19_,
         u4_sll_454_ML_int_2__20_, u4_sll_454_ML_int_2__21_,
         u4_sll_454_ML_int_2__22_, u4_sll_454_ML_int_2__23_,
         u4_sll_454_ML_int_2__24_, u4_sll_454_ML_int_2__25_,
         u4_sll_454_ML_int_2__26_, u4_sll_454_ML_int_2__27_,
         u4_sll_454_ML_int_2__28_, u4_sll_454_ML_int_2__29_,
         u4_sll_454_ML_int_2__30_, u4_sll_454_ML_int_2__31_,
         u4_sll_454_ML_int_2__32_, u4_sll_454_ML_int_2__33_,
         u4_sll_454_ML_int_2__34_, u4_sll_454_ML_int_2__35_,
         u4_sll_454_ML_int_2__36_, u4_sll_454_ML_int_2__37_,
         u4_sll_454_ML_int_2__38_, u4_sll_454_ML_int_2__39_,
         u4_sll_454_ML_int_2__40_, u4_sll_454_ML_int_2__41_,
         u4_sll_454_ML_int_2__42_, u4_sll_454_ML_int_2__43_,
         u4_sll_454_ML_int_2__44_, u4_sll_454_ML_int_2__45_,
         u4_sll_454_ML_int_2__46_, u4_sll_454_ML_int_2__47_,
         u4_sll_454_ML_int_2__48_, u4_sll_454_ML_int_2__49_,
         u4_sll_454_ML_int_2__50_, u4_sll_454_ML_int_2__51_,
         u4_sll_454_ML_int_2__52_, u4_sll_454_ML_int_2__53_,
         u4_sll_454_ML_int_2__54_, u4_sll_454_ML_int_2__55_,
         u4_sll_454_ML_int_2__56_, u4_sll_454_ML_int_2__57_,
         u4_sll_454_ML_int_2__58_, u4_sll_454_ML_int_2__59_,
         u4_sll_454_ML_int_2__60_, u4_sll_454_ML_int_2__61_,
         u4_sll_454_ML_int_2__62_, u4_sll_454_ML_int_2__63_,
         u4_sll_454_ML_int_2__64_, u4_sll_454_ML_int_2__65_,
         u4_sll_454_ML_int_2__66_, u4_sll_454_ML_int_2__67_,
         u4_sll_454_ML_int_2__68_, u4_sll_454_ML_int_2__69_,
         u4_sll_454_ML_int_2__70_, u4_sll_454_ML_int_2__71_,
         u4_sll_454_ML_int_2__72_, u4_sll_454_ML_int_2__73_,
         u4_sll_454_ML_int_2__74_, u4_sll_454_ML_int_2__75_,
         u4_sll_454_ML_int_2__76_, u4_sll_454_ML_int_2__77_,
         u4_sll_454_ML_int_2__78_, u4_sll_454_ML_int_2__79_,
         u4_sll_454_ML_int_2__80_, u4_sll_454_ML_int_2__81_,
         u4_sll_454_ML_int_2__82_, u4_sll_454_ML_int_2__83_,
         u4_sll_454_ML_int_2__84_, u4_sll_454_ML_int_2__85_,
         u4_sll_454_ML_int_2__86_, u4_sll_454_ML_int_2__87_,
         u4_sll_454_ML_int_2__88_, u4_sll_454_ML_int_2__89_,
         u4_sll_454_ML_int_2__90_, u4_sll_454_ML_int_2__91_,
         u4_sll_454_ML_int_2__92_, u4_sll_454_ML_int_2__93_,
         u4_sll_454_ML_int_2__94_, u4_sll_454_ML_int_2__95_,
         u4_sll_454_ML_int_2__96_, u4_sll_454_ML_int_2__97_,
         u4_sll_454_ML_int_2__98_, u4_sll_454_ML_int_2__99_,
         u4_sll_454_ML_int_2__100_, u4_sll_454_ML_int_2__101_,
         u4_sll_454_ML_int_2__102_, u4_sll_454_ML_int_2__103_,
         u4_sll_454_ML_int_2__104_, u4_sll_454_ML_int_2__105_,
         u4_sll_454_ML_int_1__0_, u4_sll_454_ML_int_1__1_,
         u4_sll_454_ML_int_1__2_, u4_sll_454_ML_int_1__3_,
         u4_sll_454_ML_int_1__4_, u4_sll_454_ML_int_1__5_,
         u4_sll_454_ML_int_1__6_, u4_sll_454_ML_int_1__7_,
         u4_sll_454_ML_int_1__8_, u4_sll_454_ML_int_1__9_,
         u4_sll_454_ML_int_1__10_, u4_sll_454_ML_int_1__11_,
         u4_sll_454_ML_int_1__12_, u4_sll_454_ML_int_1__13_,
         u4_sll_454_ML_int_1__14_, u4_sll_454_ML_int_1__15_,
         u4_sll_454_ML_int_1__16_, u4_sll_454_ML_int_1__17_,
         u4_sll_454_ML_int_1__18_, u4_sll_454_ML_int_1__19_,
         u4_sll_454_ML_int_1__20_, u4_sll_454_ML_int_1__21_,
         u4_sll_454_ML_int_1__22_, u4_sll_454_ML_int_1__23_,
         u4_sll_454_ML_int_1__24_, u4_sll_454_ML_int_1__25_,
         u4_sll_454_ML_int_1__26_, u4_sll_454_ML_int_1__27_,
         u4_sll_454_ML_int_1__28_, u4_sll_454_ML_int_1__29_,
         u4_sll_454_ML_int_1__30_, u4_sll_454_ML_int_1__31_,
         u4_sll_454_ML_int_1__32_, u4_sll_454_ML_int_1__33_,
         u4_sll_454_ML_int_1__34_, u4_sll_454_ML_int_1__35_,
         u4_sll_454_ML_int_1__36_, u4_sll_454_ML_int_1__37_,
         u4_sll_454_ML_int_1__38_, u4_sll_454_ML_int_1__39_,
         u4_sll_454_ML_int_1__40_, u4_sll_454_ML_int_1__41_,
         u4_sll_454_ML_int_1__42_, u4_sll_454_ML_int_1__43_,
         u4_sll_454_ML_int_1__44_, u4_sll_454_ML_int_1__45_,
         u4_sll_454_ML_int_1__46_, u4_sll_454_ML_int_1__47_,
         u4_sll_454_ML_int_1__48_, u4_sll_454_ML_int_1__49_,
         u4_sll_454_ML_int_1__50_, u4_sll_454_ML_int_1__51_,
         u4_sll_454_ML_int_1__52_, u4_sll_454_ML_int_1__53_,
         u4_sll_454_ML_int_1__54_, u4_sll_454_ML_int_1__55_,
         u4_sll_454_ML_int_1__56_, u4_sll_454_ML_int_1__57_,
         u4_sll_454_ML_int_1__58_, u4_sll_454_ML_int_1__59_,
         u4_sll_454_ML_int_1__60_, u4_sll_454_ML_int_1__61_,
         u4_sll_454_ML_int_1__62_, u4_sll_454_ML_int_1__63_,
         u4_sll_454_ML_int_1__64_, u4_sll_454_ML_int_1__65_,
         u4_sll_454_ML_int_1__66_, u4_sll_454_ML_int_1__67_,
         u4_sll_454_ML_int_1__68_, u4_sll_454_ML_int_1__69_,
         u4_sll_454_ML_int_1__70_, u4_sll_454_ML_int_1__71_,
         u4_sll_454_ML_int_1__72_, u4_sll_454_ML_int_1__73_,
         u4_sll_454_ML_int_1__74_, u4_sll_454_ML_int_1__75_,
         u4_sll_454_ML_int_1__76_, u4_sll_454_ML_int_1__77_,
         u4_sll_454_ML_int_1__78_, u4_sll_454_ML_int_1__79_,
         u4_sll_454_ML_int_1__80_, u4_sll_454_ML_int_1__81_,
         u4_sll_454_ML_int_1__82_, u4_sll_454_ML_int_1__83_,
         u4_sll_454_ML_int_1__84_, u4_sll_454_ML_int_1__85_,
         u4_sll_454_ML_int_1__86_, u4_sll_454_ML_int_1__87_,
         u4_sll_454_ML_int_1__88_, u4_sll_454_ML_int_1__89_,
         u4_sll_454_ML_int_1__90_, u4_sll_454_ML_int_1__91_,
         u4_sll_454_ML_int_1__92_, u4_sll_454_ML_int_1__93_,
         u4_sll_454_ML_int_1__94_, u4_sll_454_ML_int_1__95_,
         u4_sll_454_ML_int_1__96_, u4_sll_454_ML_int_1__97_,
         u4_sll_454_ML_int_1__98_, u4_sll_454_ML_int_1__99_,
         u4_sll_454_ML_int_1__100_, u4_sll_454_ML_int_1__101_,
         u4_sll_454_ML_int_1__102_, u4_sll_454_ML_int_1__103_,
         u4_sll_454_ML_int_1__104_, u4_sll_454_ML_int_1__105_,
         u4_sll_454_SHMAG_0_, u4_sll_454_SHMAG_1_, u4_sll_454_SHMAG_2_,
         u4_sll_454_SHMAG_3_, u4_sll_454_SHMAG_4_, u4_sll_454_SHMAG_6_,
         u4_sll_454_temp_int_SH_5_, u4_srl_453_n879, u4_srl_453_n878,
         u4_srl_453_n877, u4_srl_453_n876, u4_srl_453_n875, u4_srl_453_n874,
         u4_srl_453_n873, u4_srl_453_n872, u4_srl_453_n871, u4_srl_453_n870,
         u4_srl_453_n869, u4_srl_453_n868, u4_srl_453_n867, u4_srl_453_n866,
         u4_srl_453_n865, u4_srl_453_n864, u4_srl_453_n863, u4_srl_453_n862,
         u4_srl_453_n861, u4_srl_453_n860, u4_srl_453_n859, u4_srl_453_n858,
         u4_srl_453_n857, u4_srl_453_n856, u4_srl_453_n855, u4_srl_453_n854,
         u4_srl_453_n853, u4_srl_453_n852, u4_srl_453_n851, u4_srl_453_n850,
         u4_srl_453_n849, u4_srl_453_n848, u4_srl_453_n847, u4_srl_453_n846,
         u4_srl_453_n845, u4_srl_453_n844, u4_srl_453_n843, u4_srl_453_n842,
         u4_srl_453_n841, u4_srl_453_n840, u4_srl_453_n839, u4_srl_453_n838,
         u4_srl_453_n837, u4_srl_453_n836, u4_srl_453_n835, u4_srl_453_n834,
         u4_srl_453_n833, u4_srl_453_n832, u4_srl_453_n831, u4_srl_453_n830,
         u4_srl_453_n829, u4_srl_453_n828, u4_srl_453_n827, u4_srl_453_n826,
         u4_srl_453_n825, u4_srl_453_n824, u4_srl_453_n823, u4_srl_453_n822,
         u4_srl_453_n821, u4_srl_453_n820, u4_srl_453_n819, u4_srl_453_n818,
         u4_srl_453_n817, u4_srl_453_n816, u4_srl_453_n815, u4_srl_453_n814,
         u4_srl_453_n813, u4_srl_453_n812, u4_srl_453_n811, u4_srl_453_n810,
         u4_srl_453_n809, u4_srl_453_n808, u4_srl_453_n807, u4_srl_453_n806,
         u4_srl_453_n805, u4_srl_453_n804, u4_srl_453_n803, u4_srl_453_n802,
         u4_srl_453_n801, u4_srl_453_n800, u4_srl_453_n799, u4_srl_453_n798,
         u4_srl_453_n797, u4_srl_453_n796, u4_srl_453_n795, u4_srl_453_n794,
         u4_srl_453_n793, u4_srl_453_n792, u4_srl_453_n791, u4_srl_453_n790,
         u4_srl_453_n789, u4_srl_453_n788, u4_srl_453_n787, u4_srl_453_n786,
         u4_srl_453_n785, u4_srl_453_n784, u4_srl_453_n783, u4_srl_453_n782,
         u4_srl_453_n781, u4_srl_453_n780, u4_srl_453_n779, u4_srl_453_n778,
         u4_srl_453_n777, u4_srl_453_n776, u4_srl_453_n775, u4_srl_453_n774,
         u4_srl_453_n773, u4_srl_453_n772, u4_srl_453_n771, u4_srl_453_n770,
         u4_srl_453_n769, u4_srl_453_n768, u4_srl_453_n767, u4_srl_453_n766,
         u4_srl_453_n765, u4_srl_453_n764, u4_srl_453_n763, u4_srl_453_n762,
         u4_srl_453_n761, u4_srl_453_n760, u4_srl_453_n759, u4_srl_453_n758,
         u4_srl_453_n757, u4_srl_453_n756, u4_srl_453_n755, u4_srl_453_n754,
         u4_srl_453_n753, u4_srl_453_n752, u4_srl_453_n751, u4_srl_453_n750,
         u4_srl_453_n749, u4_srl_453_n748, u4_srl_453_n747, u4_srl_453_n746,
         u4_srl_453_n745, u4_srl_453_n744, u4_srl_453_n743, u4_srl_453_n742,
         u4_srl_453_n741, u4_srl_453_n740, u4_srl_453_n739, u4_srl_453_n738,
         u4_srl_453_n737, u4_srl_453_n736, u4_srl_453_n735, u4_srl_453_n734,
         u4_srl_453_n733, u4_srl_453_n732, u4_srl_453_n731, u4_srl_453_n730,
         u4_srl_453_n729, u4_srl_453_n728, u4_srl_453_n727, u4_srl_453_n726,
         u4_srl_453_n725, u4_srl_453_n724, u4_srl_453_n723, u4_srl_453_n722,
         u4_srl_453_n721, u4_srl_453_n720, u4_srl_453_n719, u4_srl_453_n718,
         u4_srl_453_n717, u4_srl_453_n716, u4_srl_453_n715, u4_srl_453_n714,
         u4_srl_453_n713, u4_srl_453_n712, u4_srl_453_n711, u4_srl_453_n710,
         u4_srl_453_n709, u4_srl_453_n708, u4_srl_453_n707, u4_srl_453_n706,
         u4_srl_453_n705, u4_srl_453_n704, u4_srl_453_n703, u4_srl_453_n702,
         u4_srl_453_n701, u4_srl_453_n700, u4_srl_453_n699, u4_srl_453_n698,
         u4_srl_453_n697, u4_srl_453_n696, u4_srl_453_n695, u4_srl_453_n694,
         u4_srl_453_n693, u4_srl_453_n692, u4_srl_453_n691, u4_srl_453_n690,
         u4_srl_453_n689, u4_srl_453_n688, u4_srl_453_n687, u4_srl_453_n686,
         u4_srl_453_n685, u4_srl_453_n684, u4_srl_453_n683, u4_srl_453_n682,
         u4_srl_453_n681, u4_srl_453_n680, u4_srl_453_n679, u4_srl_453_n678,
         u4_srl_453_n677, u4_srl_453_n676, u4_srl_453_n675, u4_srl_453_n674,
         u4_srl_453_n673, u4_srl_453_n672, u4_srl_453_n671, u4_srl_453_n670,
         u4_srl_453_n669, u4_srl_453_n668, u4_srl_453_n667, u4_srl_453_n666,
         u4_srl_453_n665, u4_srl_453_n664, u4_srl_453_n663, u4_srl_453_n662,
         u4_srl_453_n661, u4_srl_453_n660, u4_srl_453_n659, u4_srl_453_n658,
         u4_srl_453_n657, u4_srl_453_n656, u4_srl_453_n655, u4_srl_453_n654,
         u4_srl_453_n653, u4_srl_453_n652, u4_srl_453_n651, u4_srl_453_n650,
         u4_srl_453_n649, u4_srl_453_n648, u4_srl_453_n647, u4_srl_453_n646,
         u4_srl_453_n645, u4_srl_453_n644, u4_srl_453_n643, u4_srl_453_n642,
         u4_srl_453_n641, u4_srl_453_n640, u4_srl_453_n639, u4_srl_453_n638,
         u4_srl_453_n637, u4_srl_453_n636, u4_srl_453_n635, u4_srl_453_n634,
         u4_srl_453_n633, u4_srl_453_n632, u4_srl_453_n631, u4_srl_453_n630,
         u4_srl_453_n629, u4_srl_453_n628, u4_srl_453_n627, u4_srl_453_n626,
         u4_srl_453_n625, u4_srl_453_n624, u4_srl_453_n623, u4_srl_453_n622,
         u4_srl_453_n621, u4_srl_453_n620, u4_srl_453_n619, u4_srl_453_n618,
         u4_srl_453_n617, u4_srl_453_n616, u4_srl_453_n615, u4_srl_453_n614,
         u4_srl_453_n613, u4_srl_453_n612, u4_srl_453_n611, u4_srl_453_n610,
         u4_srl_453_n609, u4_srl_453_n608, u4_srl_453_n607, u4_srl_453_n606,
         u4_srl_453_n605, u4_srl_453_n604, u4_srl_453_n603, u4_srl_453_n602,
         u4_srl_453_n601, u4_srl_453_n600, u4_srl_453_n599, u4_srl_453_n598,
         u4_srl_453_n597, u4_srl_453_n596, u4_srl_453_n595, u4_srl_453_n594,
         u4_srl_453_n593, u4_srl_453_n592, u4_srl_453_n591, u4_srl_453_n590,
         u4_srl_453_n589, u4_srl_453_n588, u4_srl_453_n587, u4_srl_453_n586,
         u4_srl_453_n585, u4_srl_453_n584, u4_srl_453_n583, u4_srl_453_n582,
         u4_srl_453_n581, u4_srl_453_n580, u4_srl_453_n579, u4_srl_453_n578,
         u4_srl_453_n577, u4_srl_453_n576, u4_srl_453_n575, u4_srl_453_n574,
         u4_srl_453_n573, u4_srl_453_n572, u4_srl_453_n571, u4_srl_453_n570,
         u4_srl_453_n569, u4_srl_453_n568, u4_srl_453_n567, u4_srl_453_n566,
         u4_srl_453_n565, u4_srl_453_n564, u4_srl_453_n563, u4_srl_453_n562,
         u4_srl_453_n561, u4_srl_453_n560, u4_srl_453_n559, u4_srl_453_n558,
         u4_srl_453_n557, u4_srl_453_n556, u4_srl_453_n555, u4_srl_453_n554,
         u4_srl_453_n553, u4_srl_453_n552, u4_srl_453_n551, u4_srl_453_n550,
         u4_srl_453_n549, u4_srl_453_n548, u4_srl_453_n547, u4_srl_453_n546,
         u4_srl_453_n545, u4_srl_453_n544, u4_srl_453_n543, u4_srl_453_n542,
         u4_srl_453_n541, u4_srl_453_n540, u4_srl_453_n539, u4_srl_453_n538,
         u4_srl_453_n537, u4_srl_453_n536, u4_srl_453_n535, u4_srl_453_n534,
         u4_srl_453_n533, u4_srl_453_n532, u4_srl_453_n531, u4_srl_453_n530,
         u4_srl_453_n529, u4_srl_453_n528, u4_srl_453_n527, u4_srl_453_n526,
         u4_srl_453_n525, u4_srl_453_n524, u4_srl_453_n523, u4_srl_453_n522,
         u4_srl_453_n521, u4_srl_453_n520, u4_srl_453_n519, u4_srl_453_n518,
         u4_srl_453_n517, u4_srl_453_n516, u4_srl_453_n515, u4_srl_453_n514,
         u4_srl_453_n513, u4_srl_453_n512, u4_srl_453_n511, u4_srl_453_n510,
         u4_srl_453_n509, u4_srl_453_n508, u4_srl_453_n507, u4_srl_453_n506,
         u4_srl_453_n505, u4_srl_453_n504, u4_srl_453_n503, u4_srl_453_n502,
         u4_srl_453_n501, u4_srl_453_n500, u4_srl_453_n499, u4_srl_453_n498,
         u4_srl_453_n497, u4_srl_453_n496, u4_srl_453_n495, u4_srl_453_n494,
         u4_srl_453_n493, u4_srl_453_n492, u4_srl_453_n491, u4_srl_453_n490,
         u4_srl_453_n489, u4_srl_453_n488, u4_srl_453_n487, u4_srl_453_n486,
         u4_srl_453_n485, u4_srl_453_n484, u4_srl_453_n483, u4_srl_453_n482,
         u4_srl_453_n481, u4_srl_453_n480, u4_srl_453_n479, u4_srl_453_n478,
         u4_srl_453_n477, u4_srl_453_n476, u4_srl_453_n475, u4_srl_453_n474,
         u4_srl_453_n473, u4_srl_453_n472, u4_srl_453_n471, u4_srl_453_n470,
         u4_srl_453_n469, u4_srl_453_n468, u4_srl_453_n467, u4_srl_453_n466,
         u4_srl_453_n465, u4_srl_453_n464, u4_srl_453_n463, u4_srl_453_n462,
         u4_srl_453_n461, u4_srl_453_n460, u4_srl_453_n459, u4_srl_453_n458,
         u4_srl_453_n457, u4_srl_453_n456, u4_srl_453_n455, u4_srl_453_n454,
         u4_srl_453_n453, u4_srl_453_n452, u4_srl_453_n451, u4_srl_453_n450,
         u4_srl_453_n449, u4_srl_453_n448, u4_srl_453_n447, u4_srl_453_n446,
         u4_srl_453_n445, u4_srl_453_n444, u4_srl_453_n443, u4_srl_453_n442,
         u4_srl_453_n441, u4_srl_453_n440, u4_srl_453_n439, u4_srl_453_n438,
         u4_srl_453_n437, u4_srl_453_n436, u4_srl_453_n435, u4_srl_453_n434,
         u4_srl_453_n433, u4_srl_453_n432, u4_srl_453_n431, u4_srl_453_n430,
         u4_srl_453_n429, u4_srl_453_n428, u4_srl_453_n427, u4_srl_453_n426,
         u4_srl_453_n425, u4_srl_453_n424, u4_srl_453_n423, u4_srl_453_n422,
         u4_srl_453_n421, u4_srl_453_n420, u4_srl_453_n419, u4_srl_453_n418,
         u4_srl_453_n417, u4_srl_453_n416, u4_srl_453_n415, u4_srl_453_n414,
         u4_srl_453_n413, u4_srl_453_n412, u4_srl_453_n411, u4_srl_453_n410,
         u4_srl_453_n409, u4_srl_453_n408, u4_srl_453_n407, u4_srl_453_n406,
         u4_srl_453_n405, u4_srl_453_n404, u4_srl_453_n403, u4_srl_453_n402,
         u4_srl_453_n401, u4_srl_453_n400, u4_srl_453_n399, u4_srl_453_n398,
         u4_srl_453_n397, u4_srl_453_n396, u4_srl_453_n395, u4_srl_453_n394,
         u4_srl_453_n393, u4_srl_453_n392, u4_srl_453_n391, u4_srl_453_n390,
         u4_srl_453_n389, u4_srl_453_n388, u4_srl_453_n387, u4_srl_453_n386,
         u4_srl_453_n385, u4_srl_453_n384, u4_srl_453_n383, u4_srl_453_n382,
         u4_srl_453_n381, u4_srl_453_n380, u4_srl_453_n379, u4_srl_453_n378,
         u4_srl_453_n377, u4_srl_453_n376, u4_srl_453_n375, u4_srl_453_n374,
         u4_srl_453_n373, u4_srl_453_n372, u4_srl_453_n371, u4_srl_453_n370,
         u4_srl_453_n369, u4_srl_453_n368, u4_srl_453_n367, u4_srl_453_n366,
         u4_srl_453_n365, u4_srl_453_n364, u4_srl_453_n363, u4_srl_453_n362,
         u4_srl_453_n361, u4_srl_453_n360, u4_srl_453_n359, u4_srl_453_n358,
         u4_srl_453_n357, u4_srl_453_n356, u4_srl_453_n355, u4_srl_453_n354,
         u4_srl_453_n353, u4_srl_453_n352, u4_srl_453_n351, u4_srl_453_n350,
         u4_srl_453_n349, u4_srl_453_n348, u4_srl_453_n347, u4_srl_453_n346,
         u4_srl_453_n345, u4_srl_453_n344, u4_srl_453_n343, u4_srl_453_n342,
         u4_srl_453_n341, u4_srl_453_n340, u4_srl_453_n339, u4_srl_453_n338,
         u4_srl_453_n337, u4_srl_453_n336, u4_srl_453_n335, u4_srl_453_n334,
         u4_srl_453_n333, u4_srl_453_n332, u4_srl_453_n331, u4_srl_453_n330,
         u4_srl_453_n329, u4_srl_453_n328, u4_srl_453_n327, u4_srl_453_n326,
         u4_srl_453_n325, u4_srl_453_n324, u4_srl_453_n323, u4_srl_453_n322,
         u4_srl_453_n321, u4_srl_453_n320, u4_srl_453_n319, u4_srl_453_n318,
         u4_srl_453_n317, u4_srl_453_n316, u4_srl_453_n315, u4_srl_453_n314,
         u4_srl_453_n313, u4_srl_453_n312, u4_srl_453_n311, u4_srl_453_n310,
         u4_srl_453_n309, u4_srl_453_n308, u4_srl_453_n307, u4_srl_453_n306,
         u4_srl_453_n305, u4_srl_453_n304, u4_srl_453_n303, u4_srl_453_n302,
         u4_srl_453_n301, u4_srl_453_n300, u4_srl_453_n299, u4_srl_453_n298,
         u4_srl_453_n297, u4_srl_453_n296, u4_srl_453_n295, u4_srl_453_n294,
         u4_srl_453_n293, u4_srl_453_n292, u4_srl_453_n291, u4_srl_453_n290,
         u4_srl_453_n289, u4_srl_453_n288, u4_srl_453_n287, u4_srl_453_n286,
         u4_srl_453_n285, u4_srl_453_n284, u4_srl_453_n283, u4_srl_453_n282,
         u4_srl_453_n281, u4_srl_453_n280, u4_srl_453_n279, u4_srl_453_n278,
         u4_srl_453_n277, u4_srl_453_n276, u4_srl_453_n275, u4_srl_453_n274,
         u4_srl_453_n273, u4_srl_453_n272, u4_srl_453_n271, u4_srl_453_n270,
         u4_srl_453_n269, u4_srl_453_n268, u4_srl_453_n267, u4_srl_453_n266,
         u4_srl_453_n265, u4_srl_453_n264, u4_srl_453_n263, u4_srl_453_n262,
         u4_srl_453_n261, u4_srl_453_n260, u4_srl_453_n259, u4_srl_453_n258,
         u4_srl_453_n257, u4_srl_453_n256, u4_srl_453_n255, u4_srl_453_n254,
         u4_srl_453_n253, u4_srl_453_n252, u4_srl_453_n251, u4_srl_453_n250,
         u4_srl_453_n249, u4_srl_453_n248, u4_srl_453_n247, u4_srl_453_n246,
         u4_srl_453_n245, u4_srl_453_n244, u4_srl_453_n243, u4_srl_453_n242,
         u4_srl_453_n241, u4_srl_453_n240, u4_srl_453_n239, u4_srl_453_n238,
         u4_srl_453_n237, u4_srl_453_n236, u4_srl_453_n235, u4_srl_453_n234,
         u4_srl_453_n233, u4_srl_453_n232, u4_srl_453_n231, u4_srl_453_n230,
         u4_srl_453_n229, u4_srl_453_n228, u4_srl_453_n227, u4_srl_453_n226,
         u4_srl_453_n225, u4_srl_453_n224, u4_srl_453_n223, u4_srl_453_n222,
         u4_srl_453_n221, u4_srl_453_n220, u4_srl_453_n219, u4_srl_453_n218,
         u4_srl_453_n217, u4_srl_453_n216, u4_srl_453_n215, u4_srl_453_n214,
         u4_srl_453_n213, u4_srl_453_n212, u4_srl_453_n211, u4_srl_453_n210,
         u4_srl_453_n209, u4_srl_453_n208, u4_srl_453_n207, u4_srl_453_n206,
         u4_srl_453_n205, u4_srl_453_n204, u4_srl_453_n203, u4_srl_453_n202,
         u4_srl_453_n201, u4_srl_453_n200, u4_srl_453_n199, u4_srl_453_n198,
         u4_srl_453_n197, u4_srl_453_n196, u4_srl_453_n195, u4_srl_453_n194,
         u4_srl_453_n193, u4_srl_453_n192, u4_srl_453_n191, u4_srl_453_n190,
         u4_srl_453_n189, u4_srl_453_n188, u4_srl_453_n187, u4_srl_453_n186,
         u4_srl_453_n185, u4_srl_453_n184, u4_srl_453_n183, u4_srl_453_n182,
         u4_srl_453_n181, u4_srl_453_n180, u4_srl_453_n179, u4_srl_453_n178,
         u4_srl_453_n177, u4_srl_453_n176, u4_srl_453_n175, u4_srl_453_n174,
         u4_srl_453_n173, u4_srl_453_n172, u4_srl_453_n171, u4_srl_453_n170,
         u4_srl_453_n169, u4_srl_453_n168, u4_srl_453_n167, u4_srl_453_n166,
         u4_srl_453_n165, u4_srl_453_n164, u4_srl_453_n163, u4_srl_453_n162,
         u4_srl_453_n161, u4_srl_453_n160, u4_srl_453_n159, u4_srl_453_n158,
         u4_srl_453_n157, u4_srl_453_n156, u4_srl_453_n155, u4_srl_453_n154,
         u4_srl_453_n153, u4_srl_453_n152, u4_srl_453_n151, u4_srl_453_n150,
         u4_srl_453_n149, u4_srl_453_n148, u4_srl_453_n147, u4_srl_453_n146,
         u4_srl_453_n145, u4_srl_453_n144, u4_srl_453_n143, u4_srl_453_n142,
         u4_srl_453_n141, u4_srl_453_n140, u4_srl_453_n139, u4_srl_453_n138,
         u4_srl_453_n137, u4_srl_453_n136, u4_srl_453_n135, u4_srl_453_n134,
         u4_srl_453_n133, u4_srl_453_n132, u4_srl_453_n131, u4_srl_453_n130,
         u4_srl_453_n129, u4_srl_453_n128, u4_srl_453_n127, u4_srl_453_n126,
         u4_srl_453_n125, u4_srl_453_n124, u4_srl_453_n123, u4_srl_453_n122,
         u4_srl_453_n121, u4_srl_453_n120, u4_srl_453_n119, u4_srl_453_n118,
         u4_srl_453_n117, u4_srl_453_n116, u4_srl_453_n115, u4_srl_453_n114,
         u4_srl_453_n113, u4_srl_453_n112, u4_srl_453_n111, u4_srl_453_n110,
         u4_srl_453_n109, u4_srl_453_n108, u4_srl_453_n107, u4_srl_453_n106,
         u4_srl_453_n105, u4_srl_453_n104, u4_srl_453_n103, u4_srl_453_n102,
         u4_srl_453_n101, u4_srl_453_n100, u4_srl_453_n99, u4_srl_453_n98,
         u4_srl_453_n97, u4_srl_453_n96, u4_srl_453_n95, u4_srl_453_n94,
         u4_srl_453_n93, u4_srl_453_n92, u4_srl_453_n91, u4_srl_453_n90,
         u4_srl_453_n89, u4_srl_453_n88, u4_srl_453_n87, u4_srl_453_n86,
         u4_srl_453_n85, u4_srl_453_n84, u4_srl_453_n83, u4_srl_453_n82,
         u4_srl_453_n81, u4_srl_453_n80, u4_srl_453_n79, u4_srl_453_n78,
         u4_srl_453_n77, u4_srl_453_n76, u4_srl_453_n75, u4_srl_453_n74,
         u4_srl_453_n73, u4_srl_453_n72, u4_srl_453_n71, u4_srl_453_n70,
         u4_srl_453_n69, u4_srl_453_n68, u4_srl_453_n67, u4_srl_453_n66,
         u4_srl_453_n65, u4_srl_453_n64, u4_srl_453_n63, u4_srl_453_n62,
         u4_srl_453_n61, u4_srl_453_n60, u4_srl_453_n59, u4_srl_453_n58,
         u4_srl_453_n57, u4_srl_453_n56, u4_srl_453_n55, u4_srl_453_n54,
         u4_srl_453_n53, u4_srl_453_n52, u4_srl_453_n51, u4_srl_453_n50,
         u4_srl_453_n49, u4_srl_453_n48, u4_srl_453_n47, u4_srl_453_n46,
         u4_srl_453_n45, u4_srl_453_n44, u4_srl_453_n43, u4_srl_453_n42,
         u4_srl_453_n41, u4_srl_453_n40, u4_srl_453_n39, u4_srl_453_n38,
         u4_srl_453_n37, u4_srl_453_n36, u4_srl_453_n35, u4_srl_453_n34,
         u4_srl_453_n33, u4_srl_453_n32, u4_srl_453_n31, u4_srl_453_n30,
         u4_srl_453_n29, u4_srl_453_n28, u4_srl_453_n27, u4_srl_453_n26,
         u4_srl_453_n25, u4_srl_453_n24, u4_srl_453_n23, u4_srl_453_n22,
         u4_srl_453_n21, u4_srl_453_n20, u4_srl_453_n19, u4_srl_453_n18,
         u4_srl_453_n17, u4_srl_453_n16, u4_srl_453_n15, u4_srl_453_n14,
         u4_srl_453_n13, u4_srl_453_n12, u4_srl_453_n11, u4_srl_453_n10,
         u4_srl_453_n9, u4_srl_453_n8, u4_srl_453_n7, u4_srl_453_n6,
         u4_srl_453_n5, u4_srl_453_n4, u4_srl_453_n3, u4_srl_453_n2,
         u4_srl_453_n1, u4_sll_482_n57, u4_sll_482_n56, u4_sll_482_n55,
         u4_sll_482_n54, u4_sll_482_n53, u4_sll_482_n52, u4_sll_482_n51,
         u4_sll_482_n50, u4_sll_482_n49, u4_sll_482_n48, u4_sll_482_n47,
         u4_sll_482_n46, u4_sll_482_n45, u4_sll_482_n44, u4_sll_482_n43,
         u4_sll_482_n42, u4_sll_482_n41, u4_sll_482_n40, u4_sll_482_n39,
         u4_sll_482_n38, u4_sll_482_n37, u4_sll_482_n36, u4_sll_482_n35,
         u4_sll_482_n34, u4_sll_482_n33, u4_sll_482_n32, u4_sll_482_n31,
         u4_sll_482_n30, u4_sll_482_n29, u4_sll_482_n28, u4_sll_482_n27,
         u4_sll_482_n26, u4_sll_482_n25, u4_sll_482_n24, u4_sll_482_n23,
         u4_sll_482_n22, u4_sll_482_n21, u4_sll_482_n20, u4_sll_482_n19,
         u4_sll_482_n18, u4_sll_482_n17, u4_sll_482_n16, u4_sll_482_n15,
         u4_sll_482_n14, u4_sll_482_n13, u4_sll_482_n12, u4_sll_482_n11,
         u4_sll_482_n10, u4_sll_482_n9, u4_sll_482_n8, u4_sll_482_n7,
         u4_sll_482_n6, u4_sll_482_n5, u4_sll_482_n4, u4_sll_482_n3,
         u4_sll_482_n2, u4_sll_482_n1, u4_sll_482_ML_int_7__107_,
         u4_sll_482_ML_int_7__108_, u4_sll_482_ML_int_7__109_,
         u4_sll_482_ML_int_7__110_, u4_sll_482_ML_int_7__111_,
         u4_sll_482_ML_int_7__112_, u4_sll_482_ML_int_7__113_,
         u4_sll_482_ML_int_7__114_, u4_sll_482_ML_int_7__115_,
         u4_sll_482_ML_int_7__116_, u4_sll_482_ML_int_7__117_,
         u4_sll_482_ML_int_6__43_, u4_sll_482_ML_int_6__44_,
         u4_sll_482_ML_int_6__45_, u4_sll_482_ML_int_6__46_,
         u4_sll_482_ML_int_6__47_, u4_sll_482_ML_int_6__48_,
         u4_sll_482_ML_int_6__49_, u4_sll_482_ML_int_6__50_,
         u4_sll_482_ML_int_6__51_, u4_sll_482_ML_int_6__52_,
         u4_sll_482_ML_int_6__53_, u4_sll_482_ML_int_6__107_,
         u4_sll_482_ML_int_6__108_, u4_sll_482_ML_int_6__109_,
         u4_sll_482_ML_int_6__110_, u4_sll_482_ML_int_6__111_,
         u4_sll_482_ML_int_6__112_, u4_sll_482_ML_int_6__113_,
         u4_sll_482_ML_int_6__114_, u4_sll_482_ML_int_6__115_,
         u4_sll_482_ML_int_6__116_, u4_sll_482_ML_int_6__117_,
         u4_sll_482_ML_int_5__11_, u4_sll_482_ML_int_5__12_,
         u4_sll_482_ML_int_5__13_, u4_sll_482_ML_int_5__14_,
         u4_sll_482_ML_int_5__15_, u4_sll_482_ML_int_5__16_,
         u4_sll_482_ML_int_5__17_, u4_sll_482_ML_int_5__18_,
         u4_sll_482_ML_int_5__19_, u4_sll_482_ML_int_5__20_,
         u4_sll_482_ML_int_5__21_, u4_sll_482_ML_int_5__43_,
         u4_sll_482_ML_int_5__44_, u4_sll_482_ML_int_5__45_,
         u4_sll_482_ML_int_5__46_, u4_sll_482_ML_int_5__47_,
         u4_sll_482_ML_int_5__48_, u4_sll_482_ML_int_5__49_,
         u4_sll_482_ML_int_5__50_, u4_sll_482_ML_int_5__51_,
         u4_sll_482_ML_int_5__52_, u4_sll_482_ML_int_5__53_,
         u4_sll_482_ML_int_5__75_, u4_sll_482_ML_int_5__76_,
         u4_sll_482_ML_int_5__77_, u4_sll_482_ML_int_5__78_,
         u4_sll_482_ML_int_5__79_, u4_sll_482_ML_int_5__80_,
         u4_sll_482_ML_int_5__81_, u4_sll_482_ML_int_5__82_,
         u4_sll_482_ML_int_5__83_, u4_sll_482_ML_int_5__84_,
         u4_sll_482_ML_int_5__85_, u4_sll_482_ML_int_5__107_,
         u4_sll_482_ML_int_5__108_, u4_sll_482_ML_int_5__109_,
         u4_sll_482_ML_int_5__110_, u4_sll_482_ML_int_5__111_,
         u4_sll_482_ML_int_5__112_, u4_sll_482_ML_int_5__113_,
         u4_sll_482_ML_int_5__114_, u4_sll_482_ML_int_5__115_,
         u4_sll_482_ML_int_5__116_, u4_sll_482_ML_int_5__117_,
         u4_sll_482_ML_int_4__0_, u4_sll_482_ML_int_4__1_,
         u4_sll_482_ML_int_4__2_, u4_sll_482_ML_int_4__3_,
         u4_sll_482_ML_int_4__4_, u4_sll_482_ML_int_4__5_,
         u4_sll_482_ML_int_4__11_, u4_sll_482_ML_int_4__12_,
         u4_sll_482_ML_int_4__13_, u4_sll_482_ML_int_4__14_,
         u4_sll_482_ML_int_4__15_, u4_sll_482_ML_int_4__16_,
         u4_sll_482_ML_int_4__17_, u4_sll_482_ML_int_4__18_,
         u4_sll_482_ML_int_4__19_, u4_sll_482_ML_int_4__20_,
         u4_sll_482_ML_int_4__21_, u4_sll_482_ML_int_4__27_,
         u4_sll_482_ML_int_4__28_, u4_sll_482_ML_int_4__29_,
         u4_sll_482_ML_int_4__30_, u4_sll_482_ML_int_4__31_,
         u4_sll_482_ML_int_4__32_, u4_sll_482_ML_int_4__33_,
         u4_sll_482_ML_int_4__34_, u4_sll_482_ML_int_4__35_,
         u4_sll_482_ML_int_4__36_, u4_sll_482_ML_int_4__37_,
         u4_sll_482_ML_int_4__43_, u4_sll_482_ML_int_4__44_,
         u4_sll_482_ML_int_4__45_, u4_sll_482_ML_int_4__46_,
         u4_sll_482_ML_int_4__47_, u4_sll_482_ML_int_4__48_,
         u4_sll_482_ML_int_4__49_, u4_sll_482_ML_int_4__50_,
         u4_sll_482_ML_int_4__51_, u4_sll_482_ML_int_4__52_,
         u4_sll_482_ML_int_4__53_, u4_sll_482_ML_int_4__59_,
         u4_sll_482_ML_int_4__60_, u4_sll_482_ML_int_4__61_,
         u4_sll_482_ML_int_4__62_, u4_sll_482_ML_int_4__63_,
         u4_sll_482_ML_int_4__64_, u4_sll_482_ML_int_4__65_,
         u4_sll_482_ML_int_4__66_, u4_sll_482_ML_int_4__67_,
         u4_sll_482_ML_int_4__68_, u4_sll_482_ML_int_4__69_,
         u4_sll_482_ML_int_4__75_, u4_sll_482_ML_int_4__76_,
         u4_sll_482_ML_int_4__77_, u4_sll_482_ML_int_4__78_,
         u4_sll_482_ML_int_4__79_, u4_sll_482_ML_int_4__80_,
         u4_sll_482_ML_int_4__81_, u4_sll_482_ML_int_4__82_,
         u4_sll_482_ML_int_4__83_, u4_sll_482_ML_int_4__84_,
         u4_sll_482_ML_int_4__85_, u4_sll_482_ML_int_4__91_,
         u4_sll_482_ML_int_4__92_, u4_sll_482_ML_int_4__93_,
         u4_sll_482_ML_int_4__94_, u4_sll_482_ML_int_4__95_,
         u4_sll_482_ML_int_4__96_, u4_sll_482_ML_int_4__97_,
         u4_sll_482_ML_int_4__98_, u4_sll_482_ML_int_4__99_,
         u4_sll_482_ML_int_4__100_, u4_sll_482_ML_int_4__101_,
         u4_sll_482_ML_int_4__107_, u4_sll_482_ML_int_4__108_,
         u4_sll_482_ML_int_4__109_, u4_sll_482_ML_int_4__110_,
         u4_sll_482_ML_int_4__111_, u4_sll_482_ML_int_4__112_,
         u4_sll_482_ML_int_4__113_, u4_sll_482_ML_int_4__114_,
         u4_sll_482_ML_int_4__115_, u4_sll_482_ML_int_4__116_,
         u4_sll_482_ML_int_4__117_, u4_sll_482_ML_int_3__4_,
         u4_sll_482_ML_int_3__5_, u4_sll_482_ML_int_3__6_,
         u4_sll_482_ML_int_3__7_, u4_sll_482_ML_int_3__8_,
         u4_sll_482_ML_int_3__9_, u4_sll_482_ML_int_3__10_,
         u4_sll_482_ML_int_3__11_, u4_sll_482_ML_int_3__12_,
         u4_sll_482_ML_int_3__13_, u4_sll_482_ML_int_3__14_,
         u4_sll_482_ML_int_3__15_, u4_sll_482_ML_int_3__16_,
         u4_sll_482_ML_int_3__17_, u4_sll_482_ML_int_3__18_,
         u4_sll_482_ML_int_3__19_, u4_sll_482_ML_int_3__20_,
         u4_sll_482_ML_int_3__21_, u4_sll_482_ML_int_3__22_,
         u4_sll_482_ML_int_3__23_, u4_sll_482_ML_int_3__24_,
         u4_sll_482_ML_int_3__25_, u4_sll_482_ML_int_3__26_,
         u4_sll_482_ML_int_3__27_, u4_sll_482_ML_int_3__28_,
         u4_sll_482_ML_int_3__29_, u4_sll_482_ML_int_3__30_,
         u4_sll_482_ML_int_3__31_, u4_sll_482_ML_int_3__32_,
         u4_sll_482_ML_int_3__33_, u4_sll_482_ML_int_3__34_,
         u4_sll_482_ML_int_3__35_, u4_sll_482_ML_int_3__36_,
         u4_sll_482_ML_int_3__37_, u4_sll_482_ML_int_3__38_,
         u4_sll_482_ML_int_3__39_, u4_sll_482_ML_int_3__40_,
         u4_sll_482_ML_int_3__41_, u4_sll_482_ML_int_3__42_,
         u4_sll_482_ML_int_3__43_, u4_sll_482_ML_int_3__44_,
         u4_sll_482_ML_int_3__45_, u4_sll_482_ML_int_3__46_,
         u4_sll_482_ML_int_3__47_, u4_sll_482_ML_int_3__48_,
         u4_sll_482_ML_int_3__49_, u4_sll_482_ML_int_3__50_,
         u4_sll_482_ML_int_3__51_, u4_sll_482_ML_int_3__52_,
         u4_sll_482_ML_int_3__53_, u4_sll_482_ML_int_3__54_,
         u4_sll_482_ML_int_3__55_, u4_sll_482_ML_int_3__56_,
         u4_sll_482_ML_int_3__57_, u4_sll_482_ML_int_3__58_,
         u4_sll_482_ML_int_3__59_, u4_sll_482_ML_int_3__60_,
         u4_sll_482_ML_int_3__61_, u4_sll_482_ML_int_3__62_,
         u4_sll_482_ML_int_3__63_, u4_sll_482_ML_int_3__64_,
         u4_sll_482_ML_int_3__65_, u4_sll_482_ML_int_3__66_,
         u4_sll_482_ML_int_3__67_, u4_sll_482_ML_int_3__68_,
         u4_sll_482_ML_int_3__69_, u4_sll_482_ML_int_3__70_,
         u4_sll_482_ML_int_3__71_, u4_sll_482_ML_int_3__72_,
         u4_sll_482_ML_int_3__73_, u4_sll_482_ML_int_3__74_,
         u4_sll_482_ML_int_3__75_, u4_sll_482_ML_int_3__76_,
         u4_sll_482_ML_int_3__77_, u4_sll_482_ML_int_3__78_,
         u4_sll_482_ML_int_3__79_, u4_sll_482_ML_int_3__80_,
         u4_sll_482_ML_int_3__81_, u4_sll_482_ML_int_3__82_,
         u4_sll_482_ML_int_3__83_, u4_sll_482_ML_int_3__84_,
         u4_sll_482_ML_int_3__85_, u4_sll_482_ML_int_3__86_,
         u4_sll_482_ML_int_3__87_, u4_sll_482_ML_int_3__88_,
         u4_sll_482_ML_int_3__89_, u4_sll_482_ML_int_3__90_,
         u4_sll_482_ML_int_3__91_, u4_sll_482_ML_int_3__92_,
         u4_sll_482_ML_int_3__93_, u4_sll_482_ML_int_3__94_,
         u4_sll_482_ML_int_3__95_, u4_sll_482_ML_int_3__96_,
         u4_sll_482_ML_int_3__97_, u4_sll_482_ML_int_3__98_,
         u4_sll_482_ML_int_3__99_, u4_sll_482_ML_int_3__100_,
         u4_sll_482_ML_int_3__101_, u4_sll_482_ML_int_3__102_,
         u4_sll_482_ML_int_3__103_, u4_sll_482_ML_int_3__104_,
         u4_sll_482_ML_int_3__105_, u4_sll_482_ML_int_3__106_,
         u4_sll_482_ML_int_3__107_, u4_sll_482_ML_int_3__108_,
         u4_sll_482_ML_int_3__109_, u4_sll_482_ML_int_3__110_,
         u4_sll_482_ML_int_3__111_, u4_sll_482_ML_int_3__112_,
         u4_sll_482_ML_int_3__113_, u4_sll_482_ML_int_3__114_,
         u4_sll_482_ML_int_3__115_, u4_sll_482_ML_int_3__116_,
         u4_sll_482_ML_int_2__2_, u4_sll_482_ML_int_2__3_,
         u4_sll_482_ML_int_2__4_, u4_sll_482_ML_int_2__5_,
         u4_sll_482_ML_int_2__6_, u4_sll_482_ML_int_2__7_,
         u4_sll_482_ML_int_2__8_, u4_sll_482_ML_int_2__9_,
         u4_sll_482_ML_int_2__10_, u4_sll_482_ML_int_2__11_,
         u4_sll_482_ML_int_2__12_, u4_sll_482_ML_int_2__13_,
         u4_sll_482_ML_int_2__14_, u4_sll_482_ML_int_2__15_,
         u4_sll_482_ML_int_2__16_, u4_sll_482_ML_int_2__17_,
         u4_sll_482_ML_int_2__18_, u4_sll_482_ML_int_2__19_,
         u4_sll_482_ML_int_2__20_, u4_sll_482_ML_int_2__21_,
         u4_sll_482_ML_int_2__22_, u4_sll_482_ML_int_2__23_,
         u4_sll_482_ML_int_2__24_, u4_sll_482_ML_int_2__25_,
         u4_sll_482_ML_int_2__26_, u4_sll_482_ML_int_2__27_,
         u4_sll_482_ML_int_2__28_, u4_sll_482_ML_int_2__29_,
         u4_sll_482_ML_int_2__30_, u4_sll_482_ML_int_2__31_,
         u4_sll_482_ML_int_2__32_, u4_sll_482_ML_int_2__33_,
         u4_sll_482_ML_int_2__34_, u4_sll_482_ML_int_2__35_,
         u4_sll_482_ML_int_2__36_, u4_sll_482_ML_int_2__37_,
         u4_sll_482_ML_int_2__38_, u4_sll_482_ML_int_2__39_,
         u4_sll_482_ML_int_2__40_, u4_sll_482_ML_int_2__41_,
         u4_sll_482_ML_int_2__42_, u4_sll_482_ML_int_2__43_,
         u4_sll_482_ML_int_2__44_, u4_sll_482_ML_int_2__45_,
         u4_sll_482_ML_int_2__46_, u4_sll_482_ML_int_2__47_,
         u4_sll_482_ML_int_2__48_, u4_sll_482_ML_int_2__49_,
         u4_sll_482_ML_int_2__50_, u4_sll_482_ML_int_2__51_,
         u4_sll_482_ML_int_2__52_, u4_sll_482_ML_int_2__53_,
         u4_sll_482_ML_int_2__54_, u4_sll_482_ML_int_2__55_,
         u4_sll_482_ML_int_2__56_, u4_sll_482_ML_int_2__57_,
         u4_sll_482_ML_int_2__58_, u4_sll_482_ML_int_2__59_,
         u4_sll_482_ML_int_2__60_, u4_sll_482_ML_int_2__61_,
         u4_sll_482_ML_int_2__62_, u4_sll_482_ML_int_2__63_,
         u4_sll_482_ML_int_2__64_, u4_sll_482_ML_int_2__65_,
         u4_sll_482_ML_int_2__66_, u4_sll_482_ML_int_2__67_,
         u4_sll_482_ML_int_2__68_, u4_sll_482_ML_int_2__69_,
         u4_sll_482_ML_int_2__70_, u4_sll_482_ML_int_2__71_,
         u4_sll_482_ML_int_2__72_, u4_sll_482_ML_int_2__73_,
         u4_sll_482_ML_int_2__74_, u4_sll_482_ML_int_2__75_,
         u4_sll_482_ML_int_2__76_, u4_sll_482_ML_int_2__77_,
         u4_sll_482_ML_int_2__78_, u4_sll_482_ML_int_2__79_,
         u4_sll_482_ML_int_2__80_, u4_sll_482_ML_int_2__81_,
         u4_sll_482_ML_int_2__82_, u4_sll_482_ML_int_2__83_,
         u4_sll_482_ML_int_2__84_, u4_sll_482_ML_int_2__85_,
         u4_sll_482_ML_int_2__86_, u4_sll_482_ML_int_2__87_,
         u4_sll_482_ML_int_2__88_, u4_sll_482_ML_int_2__89_,
         u4_sll_482_ML_int_2__90_, u4_sll_482_ML_int_2__91_,
         u4_sll_482_ML_int_2__92_, u4_sll_482_ML_int_2__93_,
         u4_sll_482_ML_int_2__94_, u4_sll_482_ML_int_2__95_,
         u4_sll_482_ML_int_2__96_, u4_sll_482_ML_int_2__97_,
         u4_sll_482_ML_int_2__98_, u4_sll_482_ML_int_2__99_,
         u4_sll_482_ML_int_2__100_, u4_sll_482_ML_int_2__101_,
         u4_sll_482_ML_int_2__102_, u4_sll_482_ML_int_2__103_,
         u4_sll_482_ML_int_2__104_, u4_sll_482_ML_int_2__105_,
         u4_sll_482_ML_int_2__106_, u4_sll_482_ML_int_2__107_,
         u4_sll_482_ML_int_2__108_, u4_sll_482_ML_int_2__109_,
         u4_sll_482_ML_int_2__110_, u4_sll_482_ML_int_2__111_,
         u4_sll_482_ML_int_2__112_, u4_sll_482_ML_int_2__113_,
         u4_sll_482_ML_int_2__114_, u4_sll_482_ML_int_1__0_,
         u4_sll_482_ML_int_1__1_, u4_sll_482_ML_int_1__2_,
         u4_sll_482_ML_int_1__3_, u4_sll_482_ML_int_1__4_,
         u4_sll_482_ML_int_1__5_, u4_sll_482_ML_int_1__6_,
         u4_sll_482_ML_int_1__7_, u4_sll_482_ML_int_1__8_,
         u4_sll_482_ML_int_1__9_, u4_sll_482_ML_int_1__10_,
         u4_sll_482_ML_int_1__11_, u4_sll_482_ML_int_1__12_,
         u4_sll_482_ML_int_1__13_, u4_sll_482_ML_int_1__14_,
         u4_sll_482_ML_int_1__15_, u4_sll_482_ML_int_1__16_,
         u4_sll_482_ML_int_1__17_, u4_sll_482_ML_int_1__18_,
         u4_sll_482_ML_int_1__19_, u4_sll_482_ML_int_1__20_,
         u4_sll_482_ML_int_1__21_, u4_sll_482_ML_int_1__22_,
         u4_sll_482_ML_int_1__23_, u4_sll_482_ML_int_1__24_,
         u4_sll_482_ML_int_1__25_, u4_sll_482_ML_int_1__26_,
         u4_sll_482_ML_int_1__27_, u4_sll_482_ML_int_1__28_,
         u4_sll_482_ML_int_1__29_, u4_sll_482_ML_int_1__30_,
         u4_sll_482_ML_int_1__31_, u4_sll_482_ML_int_1__32_,
         u4_sll_482_ML_int_1__33_, u4_sll_482_ML_int_1__34_,
         u4_sll_482_ML_int_1__35_, u4_sll_482_ML_int_1__36_,
         u4_sll_482_ML_int_1__37_, u4_sll_482_ML_int_1__38_,
         u4_sll_482_ML_int_1__39_, u4_sll_482_ML_int_1__40_,
         u4_sll_482_ML_int_1__41_, u4_sll_482_ML_int_1__42_,
         u4_sll_482_ML_int_1__43_, u4_sll_482_ML_int_1__44_,
         u4_sll_482_ML_int_1__45_, u4_sll_482_ML_int_1__46_,
         u4_sll_482_ML_int_1__47_, u4_sll_482_ML_int_1__48_,
         u4_sll_482_ML_int_1__49_, u4_sll_482_ML_int_1__50_,
         u4_sll_482_ML_int_1__51_, u4_sll_482_ML_int_1__52_,
         u4_sll_482_ML_int_1__53_, u4_sll_482_ML_int_1__54_,
         u4_sll_482_ML_int_1__55_, u4_sll_482_ML_int_1__56_,
         u4_sll_482_ML_int_1__57_, u4_sll_482_ML_int_1__58_,
         u4_sll_482_ML_int_1__59_, u4_sll_482_ML_int_1__60_,
         u4_sll_482_ML_int_1__61_, u4_sll_482_ML_int_1__62_,
         u4_sll_482_ML_int_1__63_, u4_sll_482_ML_int_1__64_,
         u4_sll_482_ML_int_1__65_, u4_sll_482_ML_int_1__66_,
         u4_sll_482_ML_int_1__67_, u4_sll_482_ML_int_1__68_,
         u4_sll_482_ML_int_1__69_, u4_sll_482_ML_int_1__70_,
         u4_sll_482_ML_int_1__71_, u4_sll_482_ML_int_1__72_,
         u4_sll_482_ML_int_1__73_, u4_sll_482_ML_int_1__74_,
         u4_sll_482_ML_int_1__75_, u4_sll_482_ML_int_1__76_,
         u4_sll_482_ML_int_1__77_, u4_sll_482_ML_int_1__78_,
         u4_sll_482_ML_int_1__79_, u4_sll_482_ML_int_1__80_,
         u4_sll_482_ML_int_1__81_, u4_sll_482_ML_int_1__82_,
         u4_sll_482_ML_int_1__83_, u4_sll_482_ML_int_1__84_,
         u4_sll_482_ML_int_1__85_, u4_sll_482_ML_int_1__86_,
         u4_sll_482_ML_int_1__87_, u4_sll_482_ML_int_1__88_,
         u4_sll_482_ML_int_1__89_, u4_sll_482_ML_int_1__90_,
         u4_sll_482_ML_int_1__91_, u4_sll_482_ML_int_1__92_,
         u4_sll_482_ML_int_1__93_, u4_sll_482_ML_int_1__94_,
         u4_sll_482_ML_int_1__95_, u4_sll_482_ML_int_1__96_,
         u4_sll_482_ML_int_1__97_, u4_sll_482_ML_int_1__98_,
         u4_sll_482_ML_int_1__99_, u4_sll_482_ML_int_1__100_,
         u4_sll_482_ML_int_1__101_, u4_sll_482_ML_int_1__102_,
         u4_sll_482_ML_int_1__103_, u4_sll_482_ML_int_1__104_,
         u4_sll_482_ML_int_1__105_, u4_sll_482_ML_int_1__106_,
         u4_sll_482_ML_int_1__107_, u4_sll_482_ML_int_1__108_,
         u4_sll_482_ML_int_1__109_, u4_sll_482_ML_int_1__110_,
         u4_sll_482_ML_int_1__111_, u4_sll_482_ML_int_1__112_,
         u4_sll_482_ML_int_1__113_, u4_sll_482_MR_int_1__113_,
         u4_sll_482_temp_int_SH_0_, u4_sll_482_temp_int_SH_3_,
         u4_sll_482_temp_int_SH_4_, u4_sub_470_n16, u4_sub_470_n15,
         u4_sub_470_n14, u4_sub_470_n13, u4_sub_470_n12, u4_sub_470_n11,
         u4_sub_470_n10, u4_sub_470_n9, u4_sub_470_n8, u4_sub_470_n7,
         u4_sub_470_n6, u4_sub_470_n5, u4_sub_470_n4, u4_sub_470_n3,
         u4_sub_470_n2, u4_sub_470_n1, u4_sub_470_carry_1_,
         u4_sub_470_carry_2_, u4_sub_470_carry_3_, u4_sub_470_carry_4_,
         u4_sub_470_carry_5_, u4_sub_470_carry_6_, u4_sub_470_carry_7_,
         u4_sub_470_carry_8_, u4_sub_470_carry_9_, u4_sub_470_carry_10_,
         u4_sub_470_carry_11_, u4_sub_496_n14, u4_sub_496_n13, u4_sub_496_n12,
         u4_sub_496_n11, u4_sub_496_n10, u4_sub_496_n9, u4_sub_496_n8,
         u4_sub_496_n7, u4_sub_496_n6, u4_sub_496_n5, u4_sub_496_n4,
         u4_sub_496_n3, u4_sub_496_n2, u4_sub_496_n1, u4_sub_496_carry_1_,
         u4_sub_496_carry_2_, u4_sub_496_carry_3_, u4_sub_496_carry_4_,
         u4_sub_496_carry_5_, u4_sub_496_carry_6_, u4_sub_496_carry_7_,
         u4_sub_496_carry_8_, u4_sub_496_carry_9_, u4_sub_496_carry_10_,
         u4_add_489_n5, u4_add_489_n3, u4_add_489_carry_2_,
         u4_add_489_carry_3_, u4_add_489_carry_4_, u4_add_489_carry_5_,
         u4_add_494_n6, u4_add_494_n5, u4_add_494_n4, u4_add_494_carry_2_,
         u4_add_494_carry_3_, u4_add_494_carry_4_, u4_add_494_carry_5_,
         u4_add_494_carry_6_, u4_add_494_carry_7_, u4_add_494_carry_8_,
         u3_sub_63_n58, u3_sub_63_n57, u3_sub_63_n56, u3_sub_63_n55,
         u3_sub_63_n54, u3_sub_63_n53, u3_sub_63_n52, u3_sub_63_n51,
         u3_sub_63_n50, u3_sub_63_n49, u3_sub_63_n48, u3_sub_63_n47,
         u3_sub_63_n46, u3_sub_63_n45, u3_sub_63_n44, u3_sub_63_n43,
         u3_sub_63_n42, u3_sub_63_n41, u3_sub_63_n40, u3_sub_63_n39,
         u3_sub_63_n38, u3_sub_63_n37, u3_sub_63_n36, u3_sub_63_n35,
         u3_sub_63_n34, u3_sub_63_n33, u3_sub_63_n32, u3_sub_63_n31,
         u3_sub_63_n30, u3_sub_63_n29, u3_sub_63_n28, u3_sub_63_n27,
         u3_sub_63_n26, u3_sub_63_n25, u3_sub_63_n24, u3_sub_63_n23,
         u3_sub_63_n22, u3_sub_63_n21, u3_sub_63_n20, u3_sub_63_n19,
         u3_sub_63_n18, u3_sub_63_n17, u3_sub_63_n16, u3_sub_63_n15,
         u3_sub_63_n14, u3_sub_63_n13, u3_sub_63_n12, u3_sub_63_n11,
         u3_sub_63_n10, u3_sub_63_n9, u3_sub_63_n8, u3_sub_63_n7, u3_sub_63_n6,
         u3_sub_63_n5, u3_sub_63_n4, u3_sub_63_n3, u3_sub_63_n1, u3_add_63_n2,
         u2_add_115_n2, u2_sub_115_n13, u2_sub_115_n12, u2_sub_115_n11,
         u2_sub_115_n10, u2_sub_115_n9, u2_sub_115_n8, u2_sub_115_n7,
         u2_sub_115_n6, u2_sub_115_n5, u2_sub_115_n4, u2_sub_115_n3,
         u2_sub_115_n1, u1_gt_239_n167, u1_gt_239_n166, u1_gt_239_n165,
         u1_gt_239_n164, u1_gt_239_n163, u1_gt_239_n162, u1_gt_239_n161,
         u1_gt_239_n160, u1_gt_239_n159, u1_gt_239_n158, u1_gt_239_n157,
         u1_gt_239_n156, u1_gt_239_n155, u1_gt_239_n154, u1_gt_239_n153,
         u1_gt_239_n152, u1_gt_239_n151, u1_gt_239_n150, u1_gt_239_n149,
         u1_gt_239_n148, u1_gt_239_n147, u1_gt_239_n146, u1_gt_239_n145,
         u1_gt_239_n144, u1_gt_239_n143, u1_gt_239_n142, u1_gt_239_n141,
         u1_gt_239_n140, u1_gt_239_n139, u1_gt_239_n138, u1_gt_239_n137,
         u1_gt_239_n136, u1_gt_239_n135, u1_gt_239_n134, u1_gt_239_n133,
         u1_gt_239_n132, u1_gt_239_n131, u1_gt_239_n130, u1_gt_239_n129,
         u1_gt_239_n128, u1_gt_239_n127, u1_gt_239_n126, u1_gt_239_n125,
         u1_gt_239_n124, u1_gt_239_n123, u1_gt_239_n122, u1_gt_239_n121,
         u1_gt_239_n120, u1_gt_239_n119, u1_gt_239_n118, u1_gt_239_n117,
         u1_gt_239_n116, u1_gt_239_n115, u1_gt_239_n114, u1_gt_239_n113,
         u1_gt_239_n112, u1_gt_239_n111, u1_gt_239_n110, u1_gt_239_n109,
         u1_gt_239_n108, u1_gt_239_n107, u1_gt_239_n106, u1_gt_239_n105,
         u1_gt_239_n104, u1_gt_239_n103, u1_gt_239_n102, u1_gt_239_n101,
         u1_gt_239_n100, u1_gt_239_n99, u1_gt_239_n98, u1_gt_239_n97,
         u1_gt_239_n96, u1_gt_239_n95, u1_gt_239_n94, u1_gt_239_n93,
         u1_gt_239_n92, u1_gt_239_n91, u1_gt_239_n90, u1_gt_239_n89,
         u1_gt_239_n88, u1_gt_239_n87, u1_gt_239_n86, u1_gt_239_n85,
         u1_gt_239_n84, u1_gt_239_n83, u1_gt_239_n82, u1_gt_239_n81,
         u1_gt_239_n80, u1_gt_239_n79, u1_gt_239_n78, u1_gt_239_n77,
         u1_gt_239_n76, u1_gt_239_n75, u1_gt_239_n74, u1_gt_239_n73,
         u1_gt_239_n72, u1_gt_239_n71, u1_gt_239_n70, u1_gt_239_n69,
         u1_gt_239_n68, u1_gt_239_n67, u1_gt_239_n66, u1_gt_239_n65,
         u1_gt_239_n64, u1_gt_239_n63, u1_gt_239_n62, u1_gt_239_n61,
         u1_gt_239_n60, u1_gt_239_n59, u1_gt_239_n58, u1_gt_239_n57,
         u1_gt_239_n56, u1_gt_239_n55, u1_gt_239_n54, u1_gt_239_n53,
         u1_gt_239_n52, u1_gt_239_n51, u1_gt_239_n50, u1_gt_239_n49,
         u1_gt_239_n48, u1_gt_239_n47, u1_gt_239_n46, u1_gt_239_n45,
         u1_gt_239_n44, u1_gt_239_n43, u1_gt_239_n42, u1_gt_239_n41,
         u1_gt_239_n40, u1_gt_239_n39, u1_gt_239_n38, u1_gt_239_n37,
         u1_gt_239_n36, u1_gt_239_n35, u1_gt_239_n34, u1_gt_239_n33,
         u1_gt_239_n32, u1_gt_239_n31, u1_gt_239_n30, u1_gt_239_n29,
         u1_gt_239_n28, u1_gt_239_n27, u1_gt_239_n26, u1_gt_239_n25,
         u1_gt_239_n24, u1_gt_239_n23, u1_gt_239_n22, u1_gt_239_n21,
         u1_gt_239_n20, u1_gt_239_n19, u1_gt_239_n18, u1_gt_239_n17,
         u1_gt_239_n16, u1_gt_239_n15, u1_gt_239_n14, u1_gt_239_n13,
         u1_gt_239_n12, u1_gt_239_n11, u1_gt_239_n10, u1_gt_239_n9,
         u1_gt_239_n8, u1_gt_239_n7, u1_gt_239_n6, u1_gt_239_n5, u1_gt_239_n4,
         u1_gt_239_n3, u1_gt_239_n2, u1_gt_239_n1, u1_srl_151_n360,
         u1_srl_151_n359, u1_srl_151_n358, u1_srl_151_n357, u1_srl_151_n356,
         u1_srl_151_n355, u1_srl_151_n354, u1_srl_151_n353, u1_srl_151_n352,
         u1_srl_151_n351, u1_srl_151_n350, u1_srl_151_n349, u1_srl_151_n348,
         u1_srl_151_n347, u1_srl_151_n346, u1_srl_151_n345, u1_srl_151_n344,
         u1_srl_151_n343, u1_srl_151_n342, u1_srl_151_n341, u1_srl_151_n340,
         u1_srl_151_n339, u1_srl_151_n338, u1_srl_151_n337, u1_srl_151_n336,
         u1_srl_151_n335, u1_srl_151_n334, u1_srl_151_n333, u1_srl_151_n332,
         u1_srl_151_n331, u1_srl_151_n330, u1_srl_151_n329, u1_srl_151_n328,
         u1_srl_151_n327, u1_srl_151_n326, u1_srl_151_n325, u1_srl_151_n324,
         u1_srl_151_n323, u1_srl_151_n322, u1_srl_151_n321, u1_srl_151_n320,
         u1_srl_151_n319, u1_srl_151_n318, u1_srl_151_n317, u1_srl_151_n316,
         u1_srl_151_n315, u1_srl_151_n314, u1_srl_151_n313, u1_srl_151_n312,
         u1_srl_151_n311, u1_srl_151_n310, u1_srl_151_n309, u1_srl_151_n308,
         u1_srl_151_n307, u1_srl_151_n306, u1_srl_151_n305, u1_srl_151_n304,
         u1_srl_151_n303, u1_srl_151_n302, u1_srl_151_n301, u1_srl_151_n300,
         u1_srl_151_n299, u1_srl_151_n298, u1_srl_151_n297, u1_srl_151_n296,
         u1_srl_151_n295, u1_srl_151_n294, u1_srl_151_n293, u1_srl_151_n292,
         u1_srl_151_n291, u1_srl_151_n290, u1_srl_151_n289, u1_srl_151_n288,
         u1_srl_151_n287, u1_srl_151_n286, u1_srl_151_n285, u1_srl_151_n284,
         u1_srl_151_n283, u1_srl_151_n282, u1_srl_151_n281, u1_srl_151_n280,
         u1_srl_151_n279, u1_srl_151_n278, u1_srl_151_n277, u1_srl_151_n276,
         u1_srl_151_n275, u1_srl_151_n274, u1_srl_151_n273, u1_srl_151_n272,
         u1_srl_151_n271, u1_srl_151_n270, u1_srl_151_n269, u1_srl_151_n268,
         u1_srl_151_n267, u1_srl_151_n266, u1_srl_151_n265, u1_srl_151_n264,
         u1_srl_151_n263, u1_srl_151_n262, u1_srl_151_n261, u1_srl_151_n260,
         u1_srl_151_n259, u1_srl_151_n258, u1_srl_151_n257, u1_srl_151_n256,
         u1_srl_151_n255, u1_srl_151_n254, u1_srl_151_n253, u1_srl_151_n252,
         u1_srl_151_n251, u1_srl_151_n250, u1_srl_151_n249, u1_srl_151_n248,
         u1_srl_151_n247, u1_srl_151_n246, u1_srl_151_n245, u1_srl_151_n244,
         u1_srl_151_n243, u1_srl_151_n242, u1_srl_151_n241, u1_srl_151_n240,
         u1_srl_151_n239, u1_srl_151_n238, u1_srl_151_n237, u1_srl_151_n236,
         u1_srl_151_n235, u1_srl_151_n234, u1_srl_151_n233, u1_srl_151_n232,
         u1_srl_151_n231, u1_srl_151_n230, u1_srl_151_n229, u1_srl_151_n228,
         u1_srl_151_n227, u1_srl_151_n226, u1_srl_151_n225, u1_srl_151_n224,
         u1_srl_151_n223, u1_srl_151_n222, u1_srl_151_n221, u1_srl_151_n220,
         u1_srl_151_n219, u1_srl_151_n218, u1_srl_151_n217, u1_srl_151_n216,
         u1_srl_151_n215, u1_srl_151_n214, u1_srl_151_n213, u1_srl_151_n212,
         u1_srl_151_n211, u1_srl_151_n210, u1_srl_151_n209, u1_srl_151_n208,
         u1_srl_151_n207, u1_srl_151_n206, u1_srl_151_n205, u1_srl_151_n204,
         u1_srl_151_n203, u1_srl_151_n202, u1_srl_151_n201, u1_srl_151_n200,
         u1_srl_151_n199, u1_srl_151_n198, u1_srl_151_n197, u1_srl_151_n196,
         u1_srl_151_n195, u1_srl_151_n194, u1_srl_151_n193, u1_srl_151_n192,
         u1_srl_151_n191, u1_srl_151_n190, u1_srl_151_n189, u1_srl_151_n188,
         u1_srl_151_n187, u1_srl_151_n186, u1_srl_151_n185, u1_srl_151_n184,
         u1_srl_151_n183, u1_srl_151_n182, u1_srl_151_n181, u1_srl_151_n180,
         u1_srl_151_n179, u1_srl_151_n178, u1_srl_151_n177, u1_srl_151_n176,
         u1_srl_151_n175, u1_srl_151_n174, u1_srl_151_n173, u1_srl_151_n172,
         u1_srl_151_n171, u1_srl_151_n170, u1_srl_151_n169, u1_srl_151_n168,
         u1_srl_151_n167, u1_srl_151_n166, u1_srl_151_n165, u1_srl_151_n164,
         u1_srl_151_n163, u1_srl_151_n162, u1_srl_151_n161, u1_srl_151_n160,
         u1_srl_151_n159, u1_srl_151_n158, u1_srl_151_n157, u1_srl_151_n156,
         u1_srl_151_n155, u1_srl_151_n154, u1_srl_151_n153, u1_srl_151_n152,
         u1_srl_151_n151, u1_srl_151_n150, u1_srl_151_n149, u1_srl_151_n148,
         u1_srl_151_n147, u1_srl_151_n146, u1_srl_151_n145, u1_srl_151_n144,
         u1_srl_151_n143, u1_srl_151_n142, u1_srl_151_n141, u1_srl_151_n140,
         u1_srl_151_n139, u1_srl_151_n138, u1_srl_151_n137, u1_srl_151_n136,
         u1_srl_151_n135, u1_srl_151_n134, u1_srl_151_n133, u1_srl_151_n132,
         u1_srl_151_n131, u1_srl_151_n130, u1_srl_151_n129, u1_srl_151_n128,
         u1_srl_151_n127, u1_srl_151_n126, u1_srl_151_n125, u1_srl_151_n124,
         u1_srl_151_n123, u1_srl_151_n122, u1_srl_151_n121, u1_srl_151_n120,
         u1_srl_151_n119, u1_srl_151_n118, u1_srl_151_n117, u1_srl_151_n116,
         u1_srl_151_n115, u1_srl_151_n114, u1_srl_151_n113, u1_srl_151_n112,
         u1_srl_151_n111, u1_srl_151_n110, u1_srl_151_n109, u1_srl_151_n108,
         u1_srl_151_n107, u1_srl_151_n106, u1_srl_151_n105, u1_srl_151_n104,
         u1_srl_151_n103, u1_srl_151_n102, u1_srl_151_n101, u1_srl_151_n100,
         u1_srl_151_n99, u1_srl_151_n98, u1_srl_151_n97, u1_srl_151_n96,
         u1_srl_151_n95, u1_srl_151_n94, u1_srl_151_n93, u1_srl_151_n92,
         u1_srl_151_n91, u1_srl_151_n90, u1_srl_151_n89, u1_srl_151_n88,
         u1_srl_151_n87, u1_srl_151_n86, u1_srl_151_n85, u1_srl_151_n84,
         u1_srl_151_n83, u1_srl_151_n82, u1_srl_151_n81, u1_srl_151_n80,
         u1_srl_151_n79, u1_srl_151_n78, u1_srl_151_n77, u1_srl_151_n76,
         u1_srl_151_n75, u1_srl_151_n74, u1_srl_151_n73, u1_srl_151_n72,
         u1_srl_151_n71, u1_srl_151_n70, u1_srl_151_n69, u1_srl_151_n68,
         u1_srl_151_n67, u1_srl_151_n66, u1_srl_151_n65, u1_srl_151_n64,
         u1_srl_151_n63, u1_srl_151_n62, u1_srl_151_n61, u1_srl_151_n60,
         u1_srl_151_n59, u1_srl_151_n58, u1_srl_151_n57, u1_srl_151_n56,
         u1_srl_151_n55, u1_srl_151_n54, u1_srl_151_n53, u1_srl_151_n52,
         u1_srl_151_n51, u1_srl_151_n50, u1_srl_151_n49, u1_srl_151_n48,
         u1_srl_151_n47, u1_srl_151_n46, u1_srl_151_n45, u1_srl_151_n44,
         u1_srl_151_n43, u1_srl_151_n42, u1_srl_151_n41, u1_srl_151_n40,
         u1_srl_151_n39, u1_srl_151_n38, u1_srl_151_n37, u1_srl_151_n36,
         u1_srl_151_n35, u1_srl_151_n34, u1_srl_151_n33, u1_srl_151_n32,
         u1_srl_151_n31, u1_srl_151_n30, u1_srl_151_n29, u1_srl_151_n28,
         u1_srl_151_n27, u1_srl_151_n26, u1_srl_151_n25, u1_srl_151_n24,
         u1_srl_151_n23, u1_srl_151_n22, u1_srl_151_n21, u1_srl_151_n20,
         u1_srl_151_n19, u1_srl_151_n18, u1_srl_151_n17, u1_srl_151_n16,
         u1_srl_151_n15, u1_srl_151_n14, u1_srl_151_n13, u1_srl_151_n12,
         u1_srl_151_n11, u1_srl_151_n10, u1_srl_151_n9, u1_srl_151_n8,
         u1_srl_151_n7, u1_srl_151_n6, u1_srl_151_n5, u1_srl_151_n4,
         u1_srl_151_n3, u1_srl_151_n2, u1_srl_151_n1,
         sub_1_root_u1_sub_133_aco_n12, sub_1_root_u1_sub_133_aco_n11,
         sub_1_root_u1_sub_133_aco_n10, sub_1_root_u1_sub_133_aco_n9,
         sub_1_root_u1_sub_133_aco_n8, sub_1_root_u1_sub_133_aco_n7,
         sub_1_root_u1_sub_133_aco_n6, sub_1_root_u1_sub_133_aco_n5,
         sub_1_root_u1_sub_133_aco_n4, sub_1_root_u1_sub_133_aco_n3,
         sub_1_root_u1_sub_133_aco_n2, sub_1_root_u1_sub_133_aco_n1,
         sub_436_3_n171, sub_436_3_n170, sub_436_3_n169, sub_436_3_n168,
         sub_436_3_n167, sub_436_3_n166, sub_436_3_n165, sub_436_3_n164,
         sub_436_3_n163, sub_436_3_n162, sub_436_3_n161, sub_436_3_n160,
         sub_436_3_n159, sub_436_3_n158, sub_436_3_n157, sub_436_3_n156,
         sub_436_3_n155, sub_436_3_n154, sub_436_3_n153, sub_436_3_n152,
         sub_436_3_n151, sub_436_3_n150, sub_436_3_n149, sub_436_3_n148,
         sub_436_3_n147, sub_436_3_n146, sub_436_3_n145, sub_436_3_n144,
         sub_436_3_n143, sub_436_3_n142, sub_436_3_n141, sub_436_3_n140,
         sub_436_3_n139, sub_436_3_n138, sub_436_3_n137, sub_436_3_n136,
         sub_436_3_n135, sub_436_3_n134, sub_436_3_n133, sub_436_3_n132,
         sub_436_3_n131, sub_436_3_n130, sub_436_3_n129, sub_436_3_n128,
         sub_436_3_n127, sub_436_3_n126, sub_436_3_n125, sub_436_3_n124,
         sub_436_3_n123, sub_436_3_n122, sub_436_3_n121, sub_436_3_n120,
         sub_436_3_n119, sub_436_3_n118, sub_436_3_n117, sub_436_3_n116,
         sub_436_3_n115, sub_436_3_n114, sub_436_3_n97, sub_436_3_n95,
         sub_436_3_n94, sub_436_3_n93, sub_436_3_n92, sub_436_3_n91,
         sub_436_3_n90, sub_436_3_n89, sub_436_3_n88, sub_436_3_n87,
         sub_436_3_n86, sub_436_3_n85, sub_436_3_n84, sub_436_3_n83,
         sub_436_3_n82, sub_436_3_n81, sub_436_3_n80, sub_436_3_n79,
         sub_436_3_n78, sub_436_3_n77, sub_436_3_n76, sub_436_3_n52,
         sub_436_3_n51, sub_436_3_n50, sub_436_3_n49, sub_436_3_n48,
         sub_436_3_n47, sub_436_3_n46, sub_436_3_n45, sub_436_3_n44,
         sub_436_3_n43, sub_436_3_n42, sub_436_3_n41, sub_436_3_n40,
         sub_436_3_n39, sub_436_3_n38, sub_436_3_n37, sub_436_3_n36,
         sub_436_3_n23, sub_436_3_n22, sub_436_3_n21, sub_436_3_n20,
         sub_436_3_n19, sub_436_3_n18, sub_436_3_n17, sub_436_3_n16,
         sub_436_3_n15, sub_436_3_n14, sub_436_3_n13, sub_436_3_n12,
         sub_436_3_n11, sub_436_3_n10, sub_436_3_n9, sub_436_3_n8,
         sub_436_3_n7, sub_436_3_n6, sub_436_b0_n157, sub_436_b0_n156,
         sub_436_b0_n155, sub_436_b0_n154, sub_436_b0_n153, sub_436_b0_n152,
         sub_436_b0_n151, sub_436_b0_n150, sub_436_b0_n149, sub_436_b0_n148,
         sub_436_b0_n147, sub_436_b0_n146, sub_436_b0_n145, sub_436_b0_n144,
         sub_436_b0_n143, sub_436_b0_n142, sub_436_b0_n141, sub_436_b0_n140,
         sub_436_b0_n139, sub_436_b0_n138, sub_436_b0_n137, sub_436_b0_n136,
         sub_436_b0_n135, sub_436_b0_n134, sub_436_b0_n133, sub_436_b0_n132,
         sub_436_b0_n131, sub_436_b0_n130, sub_436_b0_n129, sub_436_b0_n128,
         sub_436_b0_n127, sub_436_b0_n126, sub_436_b0_n125, sub_436_b0_n124,
         sub_436_b0_n123, sub_436_b0_n122, sub_436_b0_n121, sub_436_b0_n120,
         sub_436_b0_n119, sub_436_b0_n118, sub_436_b0_n117, sub_436_b0_n116,
         sub_436_b0_n115, sub_436_b0_n114, sub_436_b0_n113, sub_436_b0_n112,
         sub_436_b0_n111, sub_436_b0_n110, sub_436_b0_n109, sub_436_b0_n108,
         sub_436_b0_n107, sub_436_b0_n106, sub_436_b0_n105, sub_436_b0_n68,
         sub_436_b0_n67, sub_436_b0_n66, sub_436_b0_n65, sub_436_b0_n64,
         sub_436_b0_n63, sub_436_b0_n62, sub_436_b0_n61, sub_436_b0_n60,
         sub_436_b0_n59, sub_436_b0_n58, sub_436_b0_n57, sub_436_b0_n56,
         sub_436_b0_n55, sub_436_b0_n54, sub_436_b0_n53, sub_436_b0_n52,
         sub_436_b0_n51, sub_436_b0_n50, sub_436_b0_n49, sub_436_b0_n48,
         sub_436_b0_n47, sub_436_b0_n46, sub_436_b0_n45, sub_436_b0_n44,
         sub_436_b0_n34, sub_436_b0_n33, sub_436_b0_n32, sub_436_b0_n31,
         sub_436_b0_n30, sub_436_b0_n29, sub_436_b0_n28, sub_436_b0_n27,
         sub_436_b0_n26, sub_436_b0_n25, sub_436_b0_n24, sub_436_b0_n23,
         sub_436_b0_n22, sub_436_b0_n21, sub_436_b0_n20, sub_436_b0_n19,
         sub_436_b0_n18, sub_436_b0_n17, sub_436_b0_n16, sub_436_b0_n15,
         sub_436_b0_n14, sub_436_b0_n13, sub_436_b0_n12, sub_436_b0_n11,
         sub_436_b0_n10, sub_436_b0_n1, sll_386_n30, sll_386_n29, sll_386_n28,
         sll_386_n27, sll_386_n26, sll_386_n25, sll_386_n24, sll_386_n23,
         sll_386_n22, sll_386_n21, sll_386_n20, sll_386_n19, sll_386_n18,
         sll_386_n17, sll_386_n16, sll_386_n15, sll_386_n14, sll_386_n13,
         sll_386_n12, sll_386_n11, sll_386_n10, sll_386_n9, sll_386_n8,
         sll_386_n7, sll_386_n6, sll_386_n5, sll_386_n4, sll_386_n3,
         sll_386_n2, sll_386_n1, sll_386_ML_int_4__8_, sll_386_ML_int_4__9_,
         sll_386_ML_int_4__10_, sll_386_ML_int_4__11_, sll_386_ML_int_4__12_,
         sll_386_ML_int_4__13_, sll_386_ML_int_4__14_, sll_386_ML_int_4__15_,
         sll_386_ML_int_4__16_, sll_386_ML_int_4__17_, sll_386_ML_int_4__18_,
         sll_386_ML_int_4__19_, sll_386_ML_int_4__20_, sll_386_ML_int_4__21_,
         sll_386_ML_int_4__22_, sll_386_ML_int_4__23_, sll_386_ML_int_4__24_,
         sll_386_ML_int_4__25_, sll_386_ML_int_4__26_, sll_386_ML_int_4__27_,
         sll_386_ML_int_4__28_, sll_386_ML_int_4__29_, sll_386_ML_int_4__30_,
         sll_386_ML_int_4__31_, sll_386_ML_int_4__32_, sll_386_ML_int_4__33_,
         sll_386_ML_int_4__34_, sll_386_ML_int_4__35_, sll_386_ML_int_4__36_,
         sll_386_ML_int_4__37_, sll_386_ML_int_4__38_, sll_386_ML_int_4__39_,
         sll_386_ML_int_4__40_, sll_386_ML_int_4__41_, sll_386_ML_int_4__42_,
         sll_386_ML_int_4__43_, sll_386_ML_int_4__44_, sll_386_ML_int_4__45_,
         sll_386_ML_int_4__46_, sll_386_ML_int_4__47_, sll_386_ML_int_4__48_,
         sll_386_ML_int_4__49_, sll_386_ML_int_4__50_, sll_386_ML_int_4__51_,
         sll_386_ML_int_4__52_, sll_386_ML_int_3__0_, sll_386_ML_int_3__1_,
         sll_386_ML_int_3__2_, sll_386_ML_int_3__3_, sll_386_ML_int_3__4_,
         sll_386_ML_int_3__5_, sll_386_ML_int_3__6_, sll_386_ML_int_3__7_,
         sll_386_ML_int_3__8_, sll_386_ML_int_3__9_, sll_386_ML_int_3__10_,
         sll_386_ML_int_3__11_, sll_386_ML_int_3__12_, sll_386_ML_int_3__13_,
         sll_386_ML_int_3__14_, sll_386_ML_int_3__15_, sll_386_ML_int_3__16_,
         sll_386_ML_int_3__17_, sll_386_ML_int_3__18_, sll_386_ML_int_3__19_,
         sll_386_ML_int_3__20_, sll_386_ML_int_3__21_, sll_386_ML_int_3__22_,
         sll_386_ML_int_3__23_, sll_386_ML_int_3__24_, sll_386_ML_int_3__25_,
         sll_386_ML_int_3__26_, sll_386_ML_int_3__27_, sll_386_ML_int_3__28_,
         sll_386_ML_int_3__29_, sll_386_ML_int_3__30_, sll_386_ML_int_3__31_,
         sll_386_ML_int_3__32_, sll_386_ML_int_3__33_, sll_386_ML_int_3__34_,
         sll_386_ML_int_3__35_, sll_386_ML_int_3__36_, sll_386_ML_int_3__37_,
         sll_386_ML_int_3__38_, sll_386_ML_int_3__39_, sll_386_ML_int_3__40_,
         sll_386_ML_int_3__41_, sll_386_ML_int_3__42_, sll_386_ML_int_3__43_,
         sll_386_ML_int_3__44_, sll_386_ML_int_3__45_, sll_386_ML_int_3__46_,
         sll_386_ML_int_3__47_, sll_386_ML_int_3__48_, sll_386_ML_int_3__49_,
         sll_386_ML_int_3__50_, sll_386_ML_int_3__51_, sll_386_ML_int_3__52_,
         sll_386_ML_int_2__0_, sll_386_ML_int_2__1_, sll_386_ML_int_2__2_,
         sll_386_ML_int_2__3_, sll_386_ML_int_2__4_, sll_386_ML_int_2__5_,
         sll_386_ML_int_2__6_, sll_386_ML_int_2__7_, sll_386_ML_int_2__8_,
         sll_386_ML_int_2__9_, sll_386_ML_int_2__10_, sll_386_ML_int_2__11_,
         sll_386_ML_int_2__12_, sll_386_ML_int_2__13_, sll_386_ML_int_2__14_,
         sll_386_ML_int_2__15_, sll_386_ML_int_2__16_, sll_386_ML_int_2__17_,
         sll_386_ML_int_2__18_, sll_386_ML_int_2__19_, sll_386_ML_int_2__20_,
         sll_386_ML_int_2__21_, sll_386_ML_int_2__22_, sll_386_ML_int_2__23_,
         sll_386_ML_int_2__24_, sll_386_ML_int_2__25_, sll_386_ML_int_2__26_,
         sll_386_ML_int_2__27_, sll_386_ML_int_2__28_, sll_386_ML_int_2__29_,
         sll_386_ML_int_2__30_, sll_386_ML_int_2__31_, sll_386_ML_int_2__32_,
         sll_386_ML_int_2__33_, sll_386_ML_int_2__34_, sll_386_ML_int_2__35_,
         sll_386_ML_int_2__36_, sll_386_ML_int_2__37_, sll_386_ML_int_2__38_,
         sll_386_ML_int_2__39_, sll_386_ML_int_2__40_, sll_386_ML_int_2__41_,
         sll_386_ML_int_2__42_, sll_386_ML_int_2__43_, sll_386_ML_int_2__44_,
         sll_386_ML_int_2__45_, sll_386_ML_int_2__46_, sll_386_ML_int_2__47_,
         sll_386_ML_int_2__48_, sll_386_ML_int_2__49_, sll_386_ML_int_2__50_,
         sll_386_ML_int_2__51_, sll_386_ML_int_2__52_, sll_386_ML_int_1__0_,
         sll_386_ML_int_1__1_, sll_386_ML_int_1__2_, sll_386_ML_int_1__3_,
         sll_386_ML_int_1__4_, sll_386_ML_int_1__5_, sll_386_ML_int_1__6_,
         sll_386_ML_int_1__7_, sll_386_ML_int_1__8_, sll_386_ML_int_1__9_,
         sll_386_ML_int_1__10_, sll_386_ML_int_1__11_, sll_386_ML_int_1__12_,
         sll_386_ML_int_1__13_, sll_386_ML_int_1__14_, sll_386_ML_int_1__15_,
         sll_386_ML_int_1__16_, sll_386_ML_int_1__17_, sll_386_ML_int_1__18_,
         sll_386_ML_int_1__19_, sll_386_ML_int_1__20_, sll_386_ML_int_1__21_,
         sll_386_ML_int_1__22_, sll_386_ML_int_1__23_, sll_386_ML_int_1__24_,
         sll_386_ML_int_1__25_, sll_386_ML_int_1__26_, sll_386_ML_int_1__27_,
         sll_386_ML_int_1__28_, sll_386_ML_int_1__29_, sll_386_ML_int_1__30_,
         sll_386_ML_int_1__31_, sll_386_ML_int_1__32_, sll_386_ML_int_1__33_,
         sll_386_ML_int_1__34_, sll_386_ML_int_1__35_, sll_386_ML_int_1__36_,
         sll_386_ML_int_1__37_, sll_386_ML_int_1__38_, sll_386_ML_int_1__39_,
         sll_386_ML_int_1__40_, sll_386_ML_int_1__41_, sll_386_ML_int_1__42_,
         sll_386_ML_int_1__43_, sll_386_ML_int_1__44_, sll_386_ML_int_1__45_,
         sll_386_ML_int_1__46_, sll_386_ML_int_1__47_, sll_386_ML_int_1__48_,
         sll_386_ML_int_1__49_, sll_386_ML_int_1__50_, sll_386_ML_int_1__51_,
         sll_386_ML_int_1__52_, r471_n178, r471_n177, r471_n176, r471_n175,
         r471_n174, r471_n173, r471_n172, r471_n171, r471_n170, r471_n169,
         r471_n168, r471_n167, r471_n166, r471_n165, r471_n164, r471_n163,
         r471_n162, r471_n161, r471_n160, r471_n159, r471_n158, r471_n157,
         r471_n156, r471_n155, r471_n154, r471_n153, r471_n152, r471_n151,
         r471_n150, r471_n149, r471_n148, r471_n147, r471_n146, r471_n145,
         r471_n144, r471_n143, r471_n142, r471_n141, r471_n140, r471_n139,
         r471_n138, r471_n137, r471_n136, r471_n135, r471_n134, r471_n133,
         r471_n132, r471_n131, r471_n130, r471_n129, r471_n128, r471_n127,
         r471_n126, r471_n125, r471_n124, r471_n123, r471_n122, r471_n121,
         r471_n120, r471_n119, r471_n118, r471_n117, r471_n116, r471_n115,
         r471_n114, r471_n113, r471_n112, r471_n111, r471_n110, r471_n109,
         r471_n108, r471_n107, r471_n106, r471_n105, r471_n104, r471_n103,
         r471_n102, r471_n101, r471_n100, r471_n99, r471_n98, r471_n97,
         r471_n96, r471_n95, r471_n94, r471_n93, r471_n92, r471_n91, r471_n90,
         r471_n89, r471_n88, r471_n87, r471_n86, r471_n85, r471_n84, r471_n83,
         r471_n82, r471_n81, r471_n80, r471_n79, r471_n78, r471_n77, r471_n76,
         r471_n75, r471_n74, r471_n73, r471_n72, r471_n71, r471_n70, r471_n69,
         r471_n68, r471_n67, r471_n66, r471_n65, r471_n64, r471_n63, r471_n62,
         r471_n61, r471_n60, r471_n59, r471_n58, r471_n57, r471_n56, r471_n55,
         r471_n54, r471_n53, r471_n52, r471_n51, r471_n50, r471_n49, r471_n48,
         r471_n47, r471_n46, r471_n45, r471_n44, r471_n43, r471_n42, r471_n41,
         r471_n40, r471_n39, r471_n38, r471_n37, r471_n36, r471_n35, r471_n34,
         r471_n33, r471_n32, r471_n31, r471_n30, r471_n29, r471_n28, r471_n27,
         r471_n26, r471_n25, r471_n24, r471_n23, r471_n22, r471_n21, r471_n20,
         r471_n19, r471_n18, r471_n17, r471_n16, r471_n15, r471_n14, r471_n13,
         r471_n12, r471_n11, r471_n10, r471_n9, r471_n8, r471_n7, r471_n6,
         r471_n5, r471_n4, r471_n3, r471_n2, r471_n1,
         add_0_root_sub_0_root_u4_add_497_n4,
         add_0_root_sub_0_root_u4_add_497_n3,
         add_0_root_sub_0_root_u4_add_497_n2,
         add_0_root_sub_0_root_u4_add_497_carry_2_,
         add_0_root_sub_0_root_u4_add_497_carry_3_,
         add_0_root_sub_0_root_u4_add_497_carry_4_,
         add_0_root_sub_0_root_u4_add_497_carry_5_,
         add_0_root_sub_0_root_u4_add_497_carry_6_,
         add_0_root_sub_0_root_u4_add_497_carry_7_,
         add_0_root_sub_0_root_u4_add_497_carry_8_, u5_mult_82_n480,
         u5_mult_82_n479, u5_mult_82_n478, u5_mult_82_n477, u5_mult_82_n476,
         u5_mult_82_n475, u5_mult_82_n474, u5_mult_82_n473, u5_mult_82_n472,
         u5_mult_82_n471, u5_mult_82_n470, u5_mult_82_n469, u5_mult_82_n468,
         u5_mult_82_n467, u5_mult_82_n466, u5_mult_82_n465, u5_mult_82_n464,
         u5_mult_82_n463, u5_mult_82_n462, u5_mult_82_n461, u5_mult_82_n460,
         u5_mult_82_n459, u5_mult_82_n458, u5_mult_82_n457, u5_mult_82_n456,
         u5_mult_82_n455, u5_mult_82_n454, u5_mult_82_n453, u5_mult_82_n452,
         u5_mult_82_n451, u5_mult_82_n450, u5_mult_82_n449, u5_mult_82_n448,
         u5_mult_82_n447, u5_mult_82_n446, u5_mult_82_n445, u5_mult_82_n444,
         u5_mult_82_n443, u5_mult_82_n442, u5_mult_82_n441, u5_mult_82_n440,
         u5_mult_82_n439, u5_mult_82_n438, u5_mult_82_n437, u5_mult_82_n436,
         u5_mult_82_n435, u5_mult_82_n434, u5_mult_82_n433, u5_mult_82_n432,
         u5_mult_82_n431, u5_mult_82_n430, u5_mult_82_n429, u5_mult_82_n428,
         u5_mult_82_n427, u5_mult_82_n426, u5_mult_82_n425, u5_mult_82_n424,
         u5_mult_82_n423, u5_mult_82_n422, u5_mult_82_n421, u5_mult_82_n420,
         u5_mult_82_n419, u5_mult_82_n418, u5_mult_82_n417, u5_mult_82_n416,
         u5_mult_82_n415, u5_mult_82_n414, u5_mult_82_n413, u5_mult_82_n412,
         u5_mult_82_n411, u5_mult_82_n410, u5_mult_82_n409, u5_mult_82_n408,
         u5_mult_82_n407, u5_mult_82_n406, u5_mult_82_n405, u5_mult_82_n404,
         u5_mult_82_n403, u5_mult_82_n402, u5_mult_82_n401, u5_mult_82_n400,
         u5_mult_82_n399, u5_mult_82_n398, u5_mult_82_n397, u5_mult_82_n396,
         u5_mult_82_n395, u5_mult_82_n394, u5_mult_82_n393, u5_mult_82_n392,
         u5_mult_82_n391, u5_mult_82_n390, u5_mult_82_n389, u5_mult_82_n388,
         u5_mult_82_n387, u5_mult_82_n386, u5_mult_82_n385, u5_mult_82_n384,
         u5_mult_82_n383, u5_mult_82_n382, u5_mult_82_n381, u5_mult_82_n380,
         u5_mult_82_n379, u5_mult_82_n378, u5_mult_82_n377, u5_mult_82_n376,
         u5_mult_82_n375, u5_mult_82_n374, u5_mult_82_n373, u5_mult_82_n372,
         u5_mult_82_n371, u5_mult_82_n370, u5_mult_82_n369, u5_mult_82_n368,
         u5_mult_82_n367, u5_mult_82_n366, u5_mult_82_n365, u5_mult_82_n364,
         u5_mult_82_n363, u5_mult_82_n362, u5_mult_82_n361, u5_mult_82_n360,
         u5_mult_82_n359, u5_mult_82_n358, u5_mult_82_n357, u5_mult_82_n356,
         u5_mult_82_n355, u5_mult_82_n354, u5_mult_82_n353, u5_mult_82_n352,
         u5_mult_82_n351, u5_mult_82_n350, u5_mult_82_n349, u5_mult_82_n348,
         u5_mult_82_n347, u5_mult_82_n346, u5_mult_82_n345, u5_mult_82_n344,
         u5_mult_82_n343, u5_mult_82_n342, u5_mult_82_n341, u5_mult_82_n340,
         u5_mult_82_n339, u5_mult_82_n338, u5_mult_82_n337, u5_mult_82_n336,
         u5_mult_82_n335, u5_mult_82_n334, u5_mult_82_n333, u5_mult_82_n332,
         u5_mult_82_n331, u5_mult_82_n330, u5_mult_82_n329, u5_mult_82_n328,
         u5_mult_82_n327, u5_mult_82_n326, u5_mult_82_n325, u5_mult_82_n324,
         u5_mult_82_n323, u5_mult_82_n322, u5_mult_82_n321, u5_mult_82_n320,
         u5_mult_82_n319, u5_mult_82_n318, u5_mult_82_n317, u5_mult_82_n316,
         u5_mult_82_n315, u5_mult_82_n314, u5_mult_82_n313, u5_mult_82_n312,
         u5_mult_82_n311, u5_mult_82_n310, u5_mult_82_n309, u5_mult_82_n308,
         u5_mult_82_n307, u5_mult_82_n306, u5_mult_82_n305, u5_mult_82_n304,
         u5_mult_82_n303, u5_mult_82_n302, u5_mult_82_n301, u5_mult_82_n300,
         u5_mult_82_n299, u5_mult_82_n298, u5_mult_82_n297, u5_mult_82_n296,
         u5_mult_82_n295, u5_mult_82_n294, u5_mult_82_n293, u5_mult_82_n292,
         u5_mult_82_n291, u5_mult_82_n290, u5_mult_82_n289, u5_mult_82_n288,
         u5_mult_82_n287, u5_mult_82_n286, u5_mult_82_n285, u5_mult_82_n284,
         u5_mult_82_n283, u5_mult_82_n282, u5_mult_82_n281, u5_mult_82_n280,
         u5_mult_82_n279, u5_mult_82_n278, u5_mult_82_n277, u5_mult_82_n276,
         u5_mult_82_n275, u5_mult_82_n274, u5_mult_82_n273, u5_mult_82_n272,
         u5_mult_82_n271, u5_mult_82_n270, u5_mult_82_n269, u5_mult_82_n268,
         u5_mult_82_n267, u5_mult_82_n266, u5_mult_82_n265, u5_mult_82_n264,
         u5_mult_82_n263, u5_mult_82_n262, u5_mult_82_n261, u5_mult_82_n260,
         u5_mult_82_n259, u5_mult_82_n258, u5_mult_82_n257, u5_mult_82_n256,
         u5_mult_82_n255, u5_mult_82_n254, u5_mult_82_n253, u5_mult_82_n252,
         u5_mult_82_n251, u5_mult_82_n250, u5_mult_82_n249, u5_mult_82_n248,
         u5_mult_82_n247, u5_mult_82_n246, u5_mult_82_n245, u5_mult_82_n244,
         u5_mult_82_n243, u5_mult_82_n242, u5_mult_82_n241, u5_mult_82_n240,
         u5_mult_82_n239, u5_mult_82_n238, u5_mult_82_n237, u5_mult_82_n236,
         u5_mult_82_n235, u5_mult_82_n234, u5_mult_82_n233, u5_mult_82_n232,
         u5_mult_82_n231, u5_mult_82_n230, u5_mult_82_n229, u5_mult_82_n228,
         u5_mult_82_n227, u5_mult_82_n226, u5_mult_82_n225, u5_mult_82_n224,
         u5_mult_82_n223, u5_mult_82_n222, u5_mult_82_n221, u5_mult_82_n220,
         u5_mult_82_n219, u5_mult_82_n218, u5_mult_82_n217, u5_mult_82_n216,
         u5_mult_82_n215, u5_mult_82_n214, u5_mult_82_n213, u5_mult_82_n212,
         u5_mult_82_n211, u5_mult_82_n209, u5_mult_82_n208, u5_mult_82_n206,
         u5_mult_82_n205, u5_mult_82_n204, u5_mult_82_n203, u5_mult_82_n202,
         u5_mult_82_n201, u5_mult_82_n200, u5_mult_82_n199, u5_mult_82_n198,
         u5_mult_82_n197, u5_mult_82_n196, u5_mult_82_n195, u5_mult_82_n194,
         u5_mult_82_n193, u5_mult_82_n192, u5_mult_82_n191, u5_mult_82_n190,
         u5_mult_82_n189, u5_mult_82_n188, u5_mult_82_n187, u5_mult_82_n186,
         u5_mult_82_n185, u5_mult_82_n184, u5_mult_82_n183, u5_mult_82_n182,
         u5_mult_82_n181, u5_mult_82_n180, u5_mult_82_n179, u5_mult_82_n178,
         u5_mult_82_n177, u5_mult_82_n176, u5_mult_82_n175, u5_mult_82_n174,
         u5_mult_82_n173, u5_mult_82_n172, u5_mult_82_n171, u5_mult_82_n170,
         u5_mult_82_n169, u5_mult_82_n168, u5_mult_82_n167, u5_mult_82_n166,
         u5_mult_82_n165, u5_mult_82_n164, u5_mult_82_n163, u5_mult_82_n162,
         u5_mult_82_n161, u5_mult_82_n160, u5_mult_82_n159, u5_mult_82_n158,
         u5_mult_82_n157, u5_mult_82_n156, u5_mult_82_n155, u5_mult_82_n154,
         u5_mult_82_n153, u5_mult_82_n152, u5_mult_82_n151, u5_mult_82_n150,
         u5_mult_82_n149, u5_mult_82_n148, u5_mult_82_n147, u5_mult_82_n146,
         u5_mult_82_n145, u5_mult_82_n144, u5_mult_82_n143, u5_mult_82_n142,
         u5_mult_82_n141, u5_mult_82_n140, u5_mult_82_n139, u5_mult_82_n138,
         u5_mult_82_n137, u5_mult_82_n136, u5_mult_82_n135, u5_mult_82_n134,
         u5_mult_82_n133, u5_mult_82_n132, u5_mult_82_n131, u5_mult_82_n130,
         u5_mult_82_n129, u5_mult_82_n128, u5_mult_82_n127, u5_mult_82_n126,
         u5_mult_82_n125, u5_mult_82_n124, u5_mult_82_n123, u5_mult_82_n122,
         u5_mult_82_n121, u5_mult_82_n120, u5_mult_82_n119, u5_mult_82_n118,
         u5_mult_82_n117, u5_mult_82_n116, u5_mult_82_n115, u5_mult_82_n114,
         u5_mult_82_n113, u5_mult_82_n112, u5_mult_82_n111, u5_mult_82_n110,
         u5_mult_82_n109, u5_mult_82_n108, u5_mult_82_n107, u5_mult_82_n106,
         u5_mult_82_n105, u5_mult_82_n104, u5_mult_82_n103, u5_mult_82_n102,
         u5_mult_82_n101, u5_mult_82_n100, u5_mult_82_n99, u5_mult_82_n98,
         u5_mult_82_n97, u5_mult_82_n96, u5_mult_82_n95, u5_mult_82_n94,
         u5_mult_82_n93, u5_mult_82_n92, u5_mult_82_n91, u5_mult_82_n90,
         u5_mult_82_n89, u5_mult_82_n88, u5_mult_82_n87, u5_mult_82_n86,
         u5_mult_82_n85, u5_mult_82_n84, u5_mult_82_n83, u5_mult_82_n82,
         u5_mult_82_n81, u5_mult_82_n80, u5_mult_82_n79, u5_mult_82_n78,
         u5_mult_82_n77, u5_mult_82_n76, u5_mult_82_n75, u5_mult_82_n74,
         u5_mult_82_n73, u5_mult_82_n72, u5_mult_82_n71, u5_mult_82_n70,
         u5_mult_82_n69, u5_mult_82_n68, u5_mult_82_n67, u5_mult_82_n66,
         u5_mult_82_n65, u5_mult_82_n64, u5_mult_82_n63, u5_mult_82_n62,
         u5_mult_82_n61, u5_mult_82_n60, u5_mult_82_n59, u5_mult_82_n58,
         u5_mult_82_n57, u5_mult_82_n56, u5_mult_82_n55, u5_mult_82_n54,
         u5_mult_82_n53, u5_mult_82_n52, u5_mult_82_n51, u5_mult_82_n50,
         u5_mult_82_n49, u5_mult_82_n48, u5_mult_82_n47, u5_mult_82_n46,
         u5_mult_82_n45, u5_mult_82_n44, u5_mult_82_n43, u5_mult_82_n42,
         u5_mult_82_n41, u5_mult_82_n40, u5_mult_82_n39, u5_mult_82_n38,
         u5_mult_82_n37, u5_mult_82_n36, u5_mult_82_n35, u5_mult_82_n34,
         u5_mult_82_n33, u5_mult_82_n32, u5_mult_82_n31, u5_mult_82_n30,
         u5_mult_82_n29, u5_mult_82_n28, u5_mult_82_n27, u5_mult_82_n26,
         u5_mult_82_n25, u5_mult_82_n24, u5_mult_82_n23, u5_mult_82_n22,
         u5_mult_82_n21, u5_mult_82_n20, u5_mult_82_n19, u5_mult_82_n18,
         u5_mult_82_n17, u5_mult_82_n16, u5_mult_82_n15, u5_mult_82_n14,
         u5_mult_82_n13, u5_mult_82_n12, u5_mult_82_n11, u5_mult_82_n10,
         u5_mult_82_n9, u5_mult_82_n8, u5_mult_82_n7, u5_mult_82_n6,
         u5_mult_82_n5, u5_mult_82_n4, u5_mult_82_n3, u5_mult_82_SUMB_43__18_,
         u5_mult_82_SUMB_43__19_, u5_mult_82_SUMB_43__20_,
         u5_mult_82_SUMB_43__21_, u5_mult_82_SUMB_43__22_,
         u5_mult_82_SUMB_43__23_, u5_mult_82_SUMB_43__24_,
         u5_mult_82_SUMB_43__25_, u5_mult_82_SUMB_43__26_,
         u5_mult_82_SUMB_43__27_, u5_mult_82_SUMB_43__28_,
         u5_mult_82_SUMB_43__29_, u5_mult_82_SUMB_43__30_,
         u5_mult_82_SUMB_43__31_, u5_mult_82_SUMB_43__32_,
         u5_mult_82_SUMB_43__33_, u5_mult_82_SUMB_43__34_,
         u5_mult_82_SUMB_43__35_, u5_mult_82_SUMB_43__36_,
         u5_mult_82_SUMB_43__37_, u5_mult_82_SUMB_43__38_,
         u5_mult_82_SUMB_43__39_, u5_mult_82_SUMB_43__40_,
         u5_mult_82_SUMB_43__41_, u5_mult_82_SUMB_43__42_,
         u5_mult_82_SUMB_43__43_, u5_mult_82_SUMB_43__44_,
         u5_mult_82_SUMB_43__45_, u5_mult_82_SUMB_43__46_,
         u5_mult_82_SUMB_43__47_, u5_mult_82_SUMB_43__48_,
         u5_mult_82_SUMB_43__49_, u5_mult_82_SUMB_43__50_,
         u5_mult_82_SUMB_43__51_, u5_mult_82_SUMB_44__1_,
         u5_mult_82_SUMB_44__2_, u5_mult_82_SUMB_44__3_,
         u5_mult_82_SUMB_44__4_, u5_mult_82_SUMB_44__5_,
         u5_mult_82_SUMB_44__6_, u5_mult_82_SUMB_44__7_,
         u5_mult_82_SUMB_44__8_, u5_mult_82_SUMB_44__9_,
         u5_mult_82_SUMB_44__10_, u5_mult_82_SUMB_44__11_,
         u5_mult_82_SUMB_44__12_, u5_mult_82_SUMB_44__13_,
         u5_mult_82_SUMB_44__14_, u5_mult_82_SUMB_44__15_,
         u5_mult_82_SUMB_44__16_, u5_mult_82_SUMB_44__17_,
         u5_mult_82_SUMB_44__18_, u5_mult_82_SUMB_44__19_,
         u5_mult_82_SUMB_44__20_, u5_mult_82_SUMB_44__21_,
         u5_mult_82_SUMB_44__22_, u5_mult_82_SUMB_44__23_,
         u5_mult_82_SUMB_44__24_, u5_mult_82_SUMB_44__25_,
         u5_mult_82_SUMB_44__26_, u5_mult_82_SUMB_44__27_,
         u5_mult_82_SUMB_44__28_, u5_mult_82_SUMB_44__29_,
         u5_mult_82_SUMB_44__30_, u5_mult_82_SUMB_44__31_,
         u5_mult_82_SUMB_44__32_, u5_mult_82_SUMB_44__33_,
         u5_mult_82_SUMB_44__34_, u5_mult_82_SUMB_44__35_,
         u5_mult_82_SUMB_44__36_, u5_mult_82_SUMB_44__37_,
         u5_mult_82_SUMB_44__38_, u5_mult_82_SUMB_44__39_,
         u5_mult_82_SUMB_44__40_, u5_mult_82_SUMB_44__41_,
         u5_mult_82_SUMB_44__42_, u5_mult_82_SUMB_44__43_,
         u5_mult_82_SUMB_44__44_, u5_mult_82_SUMB_44__45_,
         u5_mult_82_SUMB_44__46_, u5_mult_82_SUMB_44__47_,
         u5_mult_82_SUMB_44__48_, u5_mult_82_SUMB_44__49_,
         u5_mult_82_SUMB_44__50_, u5_mult_82_SUMB_44__51_,
         u5_mult_82_SUMB_45__1_, u5_mult_82_SUMB_45__2_,
         u5_mult_82_SUMB_45__3_, u5_mult_82_SUMB_45__4_,
         u5_mult_82_SUMB_45__5_, u5_mult_82_SUMB_45__6_,
         u5_mult_82_SUMB_45__7_, u5_mult_82_SUMB_45__8_,
         u5_mult_82_SUMB_45__9_, u5_mult_82_SUMB_45__10_,
         u5_mult_82_SUMB_45__11_, u5_mult_82_SUMB_45__12_,
         u5_mult_82_SUMB_45__13_, u5_mult_82_SUMB_45__14_,
         u5_mult_82_SUMB_45__15_, u5_mult_82_SUMB_45__16_,
         u5_mult_82_SUMB_45__17_, u5_mult_82_SUMB_45__18_,
         u5_mult_82_SUMB_45__19_, u5_mult_82_SUMB_45__20_,
         u5_mult_82_SUMB_45__21_, u5_mult_82_SUMB_45__22_,
         u5_mult_82_SUMB_45__23_, u5_mult_82_SUMB_45__24_,
         u5_mult_82_SUMB_45__25_, u5_mult_82_SUMB_45__26_,
         u5_mult_82_SUMB_45__27_, u5_mult_82_SUMB_45__28_,
         u5_mult_82_SUMB_45__29_, u5_mult_82_SUMB_45__30_,
         u5_mult_82_SUMB_45__31_, u5_mult_82_SUMB_45__32_,
         u5_mult_82_SUMB_45__33_, u5_mult_82_SUMB_45__34_,
         u5_mult_82_SUMB_45__35_, u5_mult_82_SUMB_45__36_,
         u5_mult_82_SUMB_45__37_, u5_mult_82_SUMB_45__38_,
         u5_mult_82_SUMB_45__39_, u5_mult_82_SUMB_45__40_,
         u5_mult_82_SUMB_45__41_, u5_mult_82_SUMB_45__42_,
         u5_mult_82_SUMB_45__43_, u5_mult_82_SUMB_45__44_,
         u5_mult_82_SUMB_45__45_, u5_mult_82_SUMB_45__46_,
         u5_mult_82_SUMB_45__47_, u5_mult_82_SUMB_45__48_,
         u5_mult_82_SUMB_45__49_, u5_mult_82_SUMB_45__50_,
         u5_mult_82_SUMB_45__51_, u5_mult_82_SUMB_46__1_,
         u5_mult_82_SUMB_46__2_, u5_mult_82_SUMB_46__3_,
         u5_mult_82_SUMB_46__4_, u5_mult_82_SUMB_46__5_,
         u5_mult_82_SUMB_46__6_, u5_mult_82_SUMB_46__7_,
         u5_mult_82_SUMB_46__8_, u5_mult_82_SUMB_46__9_,
         u5_mult_82_SUMB_46__10_, u5_mult_82_SUMB_46__11_,
         u5_mult_82_SUMB_46__12_, u5_mult_82_SUMB_46__13_,
         u5_mult_82_SUMB_46__14_, u5_mult_82_SUMB_46__15_,
         u5_mult_82_SUMB_46__16_, u5_mult_82_SUMB_46__17_,
         u5_mult_82_SUMB_46__18_, u5_mult_82_SUMB_46__19_,
         u5_mult_82_SUMB_46__20_, u5_mult_82_SUMB_46__21_,
         u5_mult_82_SUMB_46__22_, u5_mult_82_SUMB_46__23_,
         u5_mult_82_SUMB_46__24_, u5_mult_82_SUMB_46__25_,
         u5_mult_82_SUMB_46__26_, u5_mult_82_SUMB_46__27_,
         u5_mult_82_SUMB_46__28_, u5_mult_82_SUMB_46__29_,
         u5_mult_82_SUMB_46__30_, u5_mult_82_SUMB_46__31_,
         u5_mult_82_SUMB_46__32_, u5_mult_82_SUMB_46__33_,
         u5_mult_82_SUMB_46__34_, u5_mult_82_SUMB_46__35_,
         u5_mult_82_SUMB_46__36_, u5_mult_82_SUMB_46__37_,
         u5_mult_82_SUMB_46__38_, u5_mult_82_SUMB_46__39_,
         u5_mult_82_SUMB_46__40_, u5_mult_82_SUMB_46__41_,
         u5_mult_82_SUMB_46__42_, u5_mult_82_SUMB_46__43_,
         u5_mult_82_SUMB_46__44_, u5_mult_82_SUMB_46__45_,
         u5_mult_82_SUMB_46__46_, u5_mult_82_SUMB_46__47_,
         u5_mult_82_SUMB_46__48_, u5_mult_82_SUMB_46__49_,
         u5_mult_82_SUMB_46__50_, u5_mult_82_SUMB_46__51_,
         u5_mult_82_SUMB_47__1_, u5_mult_82_SUMB_47__2_,
         u5_mult_82_SUMB_47__3_, u5_mult_82_SUMB_47__4_,
         u5_mult_82_SUMB_47__5_, u5_mult_82_SUMB_47__6_,
         u5_mult_82_SUMB_47__7_, u5_mult_82_SUMB_47__8_,
         u5_mult_82_SUMB_47__9_, u5_mult_82_SUMB_47__10_,
         u5_mult_82_SUMB_47__11_, u5_mult_82_SUMB_47__12_,
         u5_mult_82_SUMB_47__13_, u5_mult_82_SUMB_47__14_,
         u5_mult_82_SUMB_47__15_, u5_mult_82_SUMB_47__16_,
         u5_mult_82_SUMB_47__17_, u5_mult_82_SUMB_47__18_,
         u5_mult_82_SUMB_47__19_, u5_mult_82_SUMB_47__20_,
         u5_mult_82_SUMB_47__21_, u5_mult_82_SUMB_47__22_,
         u5_mult_82_SUMB_47__23_, u5_mult_82_SUMB_47__24_,
         u5_mult_82_SUMB_47__25_, u5_mult_82_SUMB_47__26_,
         u5_mult_82_SUMB_47__27_, u5_mult_82_SUMB_47__28_,
         u5_mult_82_SUMB_47__29_, u5_mult_82_SUMB_47__30_,
         u5_mult_82_SUMB_47__31_, u5_mult_82_SUMB_47__32_,
         u5_mult_82_SUMB_47__33_, u5_mult_82_SUMB_47__34_,
         u5_mult_82_SUMB_47__35_, u5_mult_82_SUMB_47__36_,
         u5_mult_82_SUMB_47__37_, u5_mult_82_SUMB_47__38_,
         u5_mult_82_SUMB_47__39_, u5_mult_82_SUMB_47__40_,
         u5_mult_82_SUMB_47__41_, u5_mult_82_SUMB_47__42_,
         u5_mult_82_SUMB_47__43_, u5_mult_82_SUMB_47__44_,
         u5_mult_82_SUMB_47__45_, u5_mult_82_SUMB_47__46_,
         u5_mult_82_SUMB_47__47_, u5_mult_82_SUMB_47__48_,
         u5_mult_82_SUMB_47__49_, u5_mult_82_SUMB_47__50_,
         u5_mult_82_SUMB_47__51_, u5_mult_82_SUMB_48__1_,
         u5_mult_82_SUMB_48__2_, u5_mult_82_SUMB_48__3_,
         u5_mult_82_SUMB_48__4_, u5_mult_82_SUMB_48__5_,
         u5_mult_82_SUMB_48__6_, u5_mult_82_SUMB_48__7_,
         u5_mult_82_SUMB_48__8_, u5_mult_82_SUMB_48__9_,
         u5_mult_82_SUMB_48__10_, u5_mult_82_SUMB_48__11_,
         u5_mult_82_SUMB_48__12_, u5_mult_82_SUMB_48__13_,
         u5_mult_82_SUMB_48__14_, u5_mult_82_SUMB_48__15_,
         u5_mult_82_SUMB_48__16_, u5_mult_82_SUMB_48__17_,
         u5_mult_82_SUMB_48__18_, u5_mult_82_SUMB_48__19_,
         u5_mult_82_SUMB_48__20_, u5_mult_82_SUMB_48__21_,
         u5_mult_82_SUMB_48__22_, u5_mult_82_SUMB_48__23_,
         u5_mult_82_SUMB_48__24_, u5_mult_82_SUMB_48__25_,
         u5_mult_82_SUMB_48__26_, u5_mult_82_SUMB_48__27_,
         u5_mult_82_SUMB_48__28_, u5_mult_82_SUMB_48__29_,
         u5_mult_82_SUMB_48__30_, u5_mult_82_SUMB_48__31_,
         u5_mult_82_SUMB_48__32_, u5_mult_82_SUMB_48__33_,
         u5_mult_82_SUMB_48__34_, u5_mult_82_SUMB_48__35_,
         u5_mult_82_SUMB_48__36_, u5_mult_82_SUMB_48__37_,
         u5_mult_82_SUMB_48__38_, u5_mult_82_SUMB_48__39_,
         u5_mult_82_SUMB_48__40_, u5_mult_82_SUMB_48__41_,
         u5_mult_82_SUMB_48__42_, u5_mult_82_SUMB_48__43_,
         u5_mult_82_SUMB_48__44_, u5_mult_82_SUMB_48__45_,
         u5_mult_82_SUMB_48__46_, u5_mult_82_SUMB_48__47_,
         u5_mult_82_SUMB_48__48_, u5_mult_82_SUMB_48__49_,
         u5_mult_82_SUMB_48__50_, u5_mult_82_SUMB_48__51_,
         u5_mult_82_SUMB_49__1_, u5_mult_82_SUMB_49__2_,
         u5_mult_82_SUMB_49__3_, u5_mult_82_SUMB_49__4_,
         u5_mult_82_SUMB_49__5_, u5_mult_82_SUMB_49__6_,
         u5_mult_82_SUMB_49__7_, u5_mult_82_SUMB_49__8_,
         u5_mult_82_SUMB_49__9_, u5_mult_82_SUMB_49__10_,
         u5_mult_82_SUMB_49__11_, u5_mult_82_SUMB_49__12_,
         u5_mult_82_SUMB_49__13_, u5_mult_82_SUMB_49__14_,
         u5_mult_82_SUMB_49__15_, u5_mult_82_SUMB_49__16_,
         u5_mult_82_SUMB_49__17_, u5_mult_82_SUMB_49__18_,
         u5_mult_82_SUMB_49__19_, u5_mult_82_SUMB_49__20_,
         u5_mult_82_SUMB_49__21_, u5_mult_82_SUMB_49__22_,
         u5_mult_82_SUMB_49__23_, u5_mult_82_SUMB_49__24_,
         u5_mult_82_SUMB_49__25_, u5_mult_82_SUMB_49__26_,
         u5_mult_82_SUMB_49__27_, u5_mult_82_SUMB_49__28_,
         u5_mult_82_SUMB_49__29_, u5_mult_82_SUMB_49__30_,
         u5_mult_82_SUMB_49__31_, u5_mult_82_SUMB_49__32_,
         u5_mult_82_SUMB_49__33_, u5_mult_82_SUMB_49__34_,
         u5_mult_82_SUMB_49__35_, u5_mult_82_SUMB_49__36_,
         u5_mult_82_SUMB_49__37_, u5_mult_82_SUMB_49__38_,
         u5_mult_82_SUMB_49__39_, u5_mult_82_SUMB_49__40_,
         u5_mult_82_SUMB_49__41_, u5_mult_82_SUMB_49__42_,
         u5_mult_82_SUMB_49__43_, u5_mult_82_SUMB_49__44_,
         u5_mult_82_SUMB_49__45_, u5_mult_82_SUMB_49__46_,
         u5_mult_82_SUMB_49__47_, u5_mult_82_SUMB_49__48_,
         u5_mult_82_SUMB_49__49_, u5_mult_82_SUMB_49__50_,
         u5_mult_82_SUMB_49__51_, u5_mult_82_SUMB_50__1_,
         u5_mult_82_SUMB_50__2_, u5_mult_82_SUMB_50__3_,
         u5_mult_82_SUMB_50__4_, u5_mult_82_SUMB_50__5_,
         u5_mult_82_SUMB_50__6_, u5_mult_82_SUMB_50__7_,
         u5_mult_82_SUMB_50__8_, u5_mult_82_SUMB_50__9_,
         u5_mult_82_SUMB_50__10_, u5_mult_82_SUMB_50__11_,
         u5_mult_82_SUMB_50__12_, u5_mult_82_SUMB_50__13_,
         u5_mult_82_SUMB_50__14_, u5_mult_82_SUMB_50__15_,
         u5_mult_82_SUMB_50__16_, u5_mult_82_SUMB_50__17_,
         u5_mult_82_SUMB_50__18_, u5_mult_82_SUMB_50__19_,
         u5_mult_82_SUMB_50__20_, u5_mult_82_SUMB_50__21_,
         u5_mult_82_SUMB_50__22_, u5_mult_82_SUMB_50__23_,
         u5_mult_82_SUMB_50__24_, u5_mult_82_SUMB_50__25_,
         u5_mult_82_SUMB_50__26_, u5_mult_82_SUMB_50__27_,
         u5_mult_82_SUMB_50__28_, u5_mult_82_SUMB_50__29_,
         u5_mult_82_SUMB_50__30_, u5_mult_82_SUMB_50__31_,
         u5_mult_82_SUMB_50__32_, u5_mult_82_SUMB_50__33_,
         u5_mult_82_SUMB_50__34_, u5_mult_82_SUMB_50__35_,
         u5_mult_82_SUMB_50__36_, u5_mult_82_SUMB_50__37_,
         u5_mult_82_SUMB_50__38_, u5_mult_82_SUMB_50__39_,
         u5_mult_82_SUMB_50__40_, u5_mult_82_SUMB_50__41_,
         u5_mult_82_SUMB_50__42_, u5_mult_82_SUMB_50__43_,
         u5_mult_82_SUMB_50__44_, u5_mult_82_SUMB_50__45_,
         u5_mult_82_SUMB_50__46_, u5_mult_82_SUMB_50__47_,
         u5_mult_82_SUMB_50__48_, u5_mult_82_SUMB_50__49_,
         u5_mult_82_SUMB_50__50_, u5_mult_82_SUMB_50__51_,
         u5_mult_82_SUMB_51__1_, u5_mult_82_SUMB_51__2_,
         u5_mult_82_SUMB_51__3_, u5_mult_82_SUMB_51__4_,
         u5_mult_82_SUMB_51__5_, u5_mult_82_SUMB_51__6_,
         u5_mult_82_SUMB_51__7_, u5_mult_82_SUMB_51__8_,
         u5_mult_82_SUMB_51__9_, u5_mult_82_SUMB_51__10_,
         u5_mult_82_SUMB_51__11_, u5_mult_82_SUMB_51__12_,
         u5_mult_82_SUMB_51__13_, u5_mult_82_SUMB_51__14_,
         u5_mult_82_SUMB_51__15_, u5_mult_82_SUMB_51__16_,
         u5_mult_82_SUMB_51__17_, u5_mult_82_SUMB_51__18_,
         u5_mult_82_SUMB_51__19_, u5_mult_82_SUMB_51__20_,
         u5_mult_82_SUMB_51__21_, u5_mult_82_SUMB_51__22_,
         u5_mult_82_SUMB_51__23_, u5_mult_82_SUMB_51__24_,
         u5_mult_82_SUMB_51__25_, u5_mult_82_SUMB_51__26_,
         u5_mult_82_SUMB_51__27_, u5_mult_82_SUMB_51__28_,
         u5_mult_82_SUMB_51__29_, u5_mult_82_SUMB_51__30_,
         u5_mult_82_SUMB_51__31_, u5_mult_82_SUMB_51__32_,
         u5_mult_82_SUMB_51__33_, u5_mult_82_SUMB_51__34_,
         u5_mult_82_SUMB_51__35_, u5_mult_82_SUMB_51__36_,
         u5_mult_82_SUMB_51__37_, u5_mult_82_SUMB_51__38_,
         u5_mult_82_SUMB_51__39_, u5_mult_82_SUMB_51__40_,
         u5_mult_82_SUMB_51__41_, u5_mult_82_SUMB_51__42_,
         u5_mult_82_SUMB_51__43_, u5_mult_82_SUMB_51__44_,
         u5_mult_82_SUMB_51__45_, u5_mult_82_SUMB_51__46_,
         u5_mult_82_SUMB_51__47_, u5_mult_82_SUMB_51__48_,
         u5_mult_82_SUMB_51__49_, u5_mult_82_SUMB_51__50_,
         u5_mult_82_SUMB_51__51_, u5_mult_82_SUMB_52__1_,
         u5_mult_82_SUMB_52__2_, u5_mult_82_SUMB_52__3_,
         u5_mult_82_SUMB_52__4_, u5_mult_82_SUMB_52__5_,
         u5_mult_82_SUMB_52__6_, u5_mult_82_SUMB_52__7_,
         u5_mult_82_SUMB_52__8_, u5_mult_82_SUMB_52__9_,
         u5_mult_82_SUMB_52__10_, u5_mult_82_SUMB_52__11_,
         u5_mult_82_SUMB_52__12_, u5_mult_82_SUMB_52__13_,
         u5_mult_82_SUMB_52__14_, u5_mult_82_SUMB_52__15_,
         u5_mult_82_SUMB_52__16_, u5_mult_82_SUMB_52__17_,
         u5_mult_82_SUMB_52__18_, u5_mult_82_SUMB_52__19_,
         u5_mult_82_SUMB_52__20_, u5_mult_82_SUMB_52__21_,
         u5_mult_82_SUMB_52__22_, u5_mult_82_SUMB_52__23_,
         u5_mult_82_SUMB_52__24_, u5_mult_82_SUMB_52__25_,
         u5_mult_82_SUMB_52__26_, u5_mult_82_SUMB_52__27_,
         u5_mult_82_SUMB_52__28_, u5_mult_82_SUMB_52__29_,
         u5_mult_82_SUMB_52__30_, u5_mult_82_SUMB_52__31_,
         u5_mult_82_SUMB_52__32_, u5_mult_82_SUMB_52__33_,
         u5_mult_82_SUMB_52__34_, u5_mult_82_SUMB_52__35_,
         u5_mult_82_SUMB_52__36_, u5_mult_82_SUMB_52__37_,
         u5_mult_82_SUMB_52__38_, u5_mult_82_SUMB_52__39_,
         u5_mult_82_SUMB_52__40_, u5_mult_82_SUMB_52__41_,
         u5_mult_82_SUMB_52__42_, u5_mult_82_SUMB_52__43_,
         u5_mult_82_SUMB_52__44_, u5_mult_82_SUMB_52__45_,
         u5_mult_82_SUMB_52__46_, u5_mult_82_SUMB_52__47_,
         u5_mult_82_SUMB_52__48_, u5_mult_82_SUMB_52__49_,
         u5_mult_82_SUMB_52__50_, u5_mult_82_SUMB_52__51_,
         u5_mult_82_CARRYB_43__18_, u5_mult_82_CARRYB_43__19_,
         u5_mult_82_CARRYB_43__20_, u5_mult_82_CARRYB_43__21_,
         u5_mult_82_CARRYB_43__22_, u5_mult_82_CARRYB_43__23_,
         u5_mult_82_CARRYB_43__24_, u5_mult_82_CARRYB_43__25_,
         u5_mult_82_CARRYB_43__26_, u5_mult_82_CARRYB_43__27_,
         u5_mult_82_CARRYB_43__28_, u5_mult_82_CARRYB_43__29_,
         u5_mult_82_CARRYB_43__30_, u5_mult_82_CARRYB_43__31_,
         u5_mult_82_CARRYB_43__32_, u5_mult_82_CARRYB_43__33_,
         u5_mult_82_CARRYB_43__34_, u5_mult_82_CARRYB_43__35_,
         u5_mult_82_CARRYB_43__36_, u5_mult_82_CARRYB_43__37_,
         u5_mult_82_CARRYB_43__38_, u5_mult_82_CARRYB_43__39_,
         u5_mult_82_CARRYB_43__40_, u5_mult_82_CARRYB_43__41_,
         u5_mult_82_CARRYB_43__42_, u5_mult_82_CARRYB_43__43_,
         u5_mult_82_CARRYB_43__44_, u5_mult_82_CARRYB_43__45_,
         u5_mult_82_CARRYB_43__46_, u5_mult_82_CARRYB_43__47_,
         u5_mult_82_CARRYB_43__48_, u5_mult_82_CARRYB_43__49_,
         u5_mult_82_CARRYB_43__50_, u5_mult_82_CARRYB_43__51_,
         u5_mult_82_CARRYB_44__0_, u5_mult_82_CARRYB_44__1_,
         u5_mult_82_CARRYB_44__2_, u5_mult_82_CARRYB_44__3_,
         u5_mult_82_CARRYB_44__4_, u5_mult_82_CARRYB_44__5_,
         u5_mult_82_CARRYB_44__6_, u5_mult_82_CARRYB_44__7_,
         u5_mult_82_CARRYB_44__8_, u5_mult_82_CARRYB_44__9_,
         u5_mult_82_CARRYB_44__10_, u5_mult_82_CARRYB_44__11_,
         u5_mult_82_CARRYB_44__12_, u5_mult_82_CARRYB_44__13_,
         u5_mult_82_CARRYB_44__14_, u5_mult_82_CARRYB_44__15_,
         u5_mult_82_CARRYB_44__16_, u5_mult_82_CARRYB_44__17_,
         u5_mult_82_CARRYB_44__18_, u5_mult_82_CARRYB_44__19_,
         u5_mult_82_CARRYB_44__20_, u5_mult_82_CARRYB_44__21_,
         u5_mult_82_CARRYB_44__22_, u5_mult_82_CARRYB_44__23_,
         u5_mult_82_CARRYB_44__24_, u5_mult_82_CARRYB_44__25_,
         u5_mult_82_CARRYB_44__26_, u5_mult_82_CARRYB_44__27_,
         u5_mult_82_CARRYB_44__28_, u5_mult_82_CARRYB_44__29_,
         u5_mult_82_CARRYB_44__30_, u5_mult_82_CARRYB_44__31_,
         u5_mult_82_CARRYB_44__32_, u5_mult_82_CARRYB_44__33_,
         u5_mult_82_CARRYB_44__34_, u5_mult_82_CARRYB_44__35_,
         u5_mult_82_CARRYB_44__36_, u5_mult_82_CARRYB_44__37_,
         u5_mult_82_CARRYB_44__38_, u5_mult_82_CARRYB_44__39_,
         u5_mult_82_CARRYB_44__40_, u5_mult_82_CARRYB_44__41_,
         u5_mult_82_CARRYB_44__42_, u5_mult_82_CARRYB_44__43_,
         u5_mult_82_CARRYB_44__44_, u5_mult_82_CARRYB_44__45_,
         u5_mult_82_CARRYB_44__46_, u5_mult_82_CARRYB_44__47_,
         u5_mult_82_CARRYB_44__48_, u5_mult_82_CARRYB_44__49_,
         u5_mult_82_CARRYB_44__50_, u5_mult_82_CARRYB_44__51_,
         u5_mult_82_CARRYB_45__0_, u5_mult_82_CARRYB_45__1_,
         u5_mult_82_CARRYB_45__2_, u5_mult_82_CARRYB_45__3_,
         u5_mult_82_CARRYB_45__4_, u5_mult_82_CARRYB_45__5_,
         u5_mult_82_CARRYB_45__6_, u5_mult_82_CARRYB_45__7_,
         u5_mult_82_CARRYB_45__8_, u5_mult_82_CARRYB_45__9_,
         u5_mult_82_CARRYB_45__10_, u5_mult_82_CARRYB_45__11_,
         u5_mult_82_CARRYB_45__12_, u5_mult_82_CARRYB_45__13_,
         u5_mult_82_CARRYB_45__14_, u5_mult_82_CARRYB_45__15_,
         u5_mult_82_CARRYB_45__16_, u5_mult_82_CARRYB_45__17_,
         u5_mult_82_CARRYB_45__18_, u5_mult_82_CARRYB_45__19_,
         u5_mult_82_CARRYB_45__20_, u5_mult_82_CARRYB_45__21_,
         u5_mult_82_CARRYB_45__22_, u5_mult_82_CARRYB_45__23_,
         u5_mult_82_CARRYB_45__24_, u5_mult_82_CARRYB_45__25_,
         u5_mult_82_CARRYB_45__26_, u5_mult_82_CARRYB_45__27_,
         u5_mult_82_CARRYB_45__28_, u5_mult_82_CARRYB_45__29_,
         u5_mult_82_CARRYB_45__30_, u5_mult_82_CARRYB_45__31_,
         u5_mult_82_CARRYB_45__32_, u5_mult_82_CARRYB_45__33_,
         u5_mult_82_CARRYB_45__34_, u5_mult_82_CARRYB_45__35_,
         u5_mult_82_CARRYB_45__36_, u5_mult_82_CARRYB_45__37_,
         u5_mult_82_CARRYB_45__38_, u5_mult_82_CARRYB_45__39_,
         u5_mult_82_CARRYB_45__40_, u5_mult_82_CARRYB_45__41_,
         u5_mult_82_CARRYB_45__42_, u5_mult_82_CARRYB_45__43_,
         u5_mult_82_CARRYB_45__44_, u5_mult_82_CARRYB_45__45_,
         u5_mult_82_CARRYB_45__46_, u5_mult_82_CARRYB_45__47_,
         u5_mult_82_CARRYB_45__48_, u5_mult_82_CARRYB_45__49_,
         u5_mult_82_CARRYB_45__50_, u5_mult_82_CARRYB_45__51_,
         u5_mult_82_CARRYB_46__0_, u5_mult_82_CARRYB_46__1_,
         u5_mult_82_CARRYB_46__2_, u5_mult_82_CARRYB_46__3_,
         u5_mult_82_CARRYB_46__4_, u5_mult_82_CARRYB_46__5_,
         u5_mult_82_CARRYB_46__6_, u5_mult_82_CARRYB_46__7_,
         u5_mult_82_CARRYB_46__8_, u5_mult_82_CARRYB_46__9_,
         u5_mult_82_CARRYB_46__10_, u5_mult_82_CARRYB_46__11_,
         u5_mult_82_CARRYB_46__12_, u5_mult_82_CARRYB_46__13_,
         u5_mult_82_CARRYB_46__14_, u5_mult_82_CARRYB_46__15_,
         u5_mult_82_CARRYB_46__16_, u5_mult_82_CARRYB_46__17_,
         u5_mult_82_CARRYB_46__18_, u5_mult_82_CARRYB_46__19_,
         u5_mult_82_CARRYB_46__20_, u5_mult_82_CARRYB_46__21_,
         u5_mult_82_CARRYB_46__22_, u5_mult_82_CARRYB_46__23_,
         u5_mult_82_CARRYB_46__24_, u5_mult_82_CARRYB_46__25_,
         u5_mult_82_CARRYB_46__26_, u5_mult_82_CARRYB_46__27_,
         u5_mult_82_CARRYB_46__28_, u5_mult_82_CARRYB_46__29_,
         u5_mult_82_CARRYB_46__30_, u5_mult_82_CARRYB_46__31_,
         u5_mult_82_CARRYB_46__32_, u5_mult_82_CARRYB_46__33_,
         u5_mult_82_CARRYB_46__34_, u5_mult_82_CARRYB_46__35_,
         u5_mult_82_CARRYB_46__36_, u5_mult_82_CARRYB_46__37_,
         u5_mult_82_CARRYB_46__38_, u5_mult_82_CARRYB_46__39_,
         u5_mult_82_CARRYB_46__40_, u5_mult_82_CARRYB_46__41_,
         u5_mult_82_CARRYB_46__42_, u5_mult_82_CARRYB_46__43_,
         u5_mult_82_CARRYB_46__44_, u5_mult_82_CARRYB_46__45_,
         u5_mult_82_CARRYB_46__46_, u5_mult_82_CARRYB_46__47_,
         u5_mult_82_CARRYB_46__48_, u5_mult_82_CARRYB_46__49_,
         u5_mult_82_CARRYB_46__50_, u5_mult_82_CARRYB_46__51_,
         u5_mult_82_CARRYB_47__0_, u5_mult_82_CARRYB_47__1_,
         u5_mult_82_CARRYB_47__2_, u5_mult_82_CARRYB_47__3_,
         u5_mult_82_CARRYB_47__4_, u5_mult_82_CARRYB_47__5_,
         u5_mult_82_CARRYB_47__6_, u5_mult_82_CARRYB_47__7_,
         u5_mult_82_CARRYB_47__8_, u5_mult_82_CARRYB_47__9_,
         u5_mult_82_CARRYB_47__10_, u5_mult_82_CARRYB_47__11_,
         u5_mult_82_CARRYB_47__12_, u5_mult_82_CARRYB_47__13_,
         u5_mult_82_CARRYB_47__14_, u5_mult_82_CARRYB_47__15_,
         u5_mult_82_CARRYB_47__16_, u5_mult_82_CARRYB_47__17_,
         u5_mult_82_CARRYB_47__18_, u5_mult_82_CARRYB_47__19_,
         u5_mult_82_CARRYB_47__20_, u5_mult_82_CARRYB_47__21_,
         u5_mult_82_CARRYB_47__22_, u5_mult_82_CARRYB_47__23_,
         u5_mult_82_CARRYB_47__24_, u5_mult_82_CARRYB_47__25_,
         u5_mult_82_CARRYB_47__26_, u5_mult_82_CARRYB_47__27_,
         u5_mult_82_CARRYB_47__28_, u5_mult_82_CARRYB_47__29_,
         u5_mult_82_CARRYB_47__30_, u5_mult_82_CARRYB_47__31_,
         u5_mult_82_CARRYB_47__32_, u5_mult_82_CARRYB_47__33_,
         u5_mult_82_CARRYB_47__34_, u5_mult_82_CARRYB_47__35_,
         u5_mult_82_CARRYB_47__36_, u5_mult_82_CARRYB_47__37_,
         u5_mult_82_CARRYB_47__38_, u5_mult_82_CARRYB_47__39_,
         u5_mult_82_CARRYB_47__40_, u5_mult_82_CARRYB_47__41_,
         u5_mult_82_CARRYB_47__42_, u5_mult_82_CARRYB_47__43_,
         u5_mult_82_CARRYB_47__44_, u5_mult_82_CARRYB_47__45_,
         u5_mult_82_CARRYB_47__46_, u5_mult_82_CARRYB_47__47_,
         u5_mult_82_CARRYB_47__48_, u5_mult_82_CARRYB_47__49_,
         u5_mult_82_CARRYB_47__50_, u5_mult_82_CARRYB_47__51_,
         u5_mult_82_CARRYB_48__0_, u5_mult_82_CARRYB_48__1_,
         u5_mult_82_CARRYB_48__2_, u5_mult_82_CARRYB_48__3_,
         u5_mult_82_CARRYB_48__4_, u5_mult_82_CARRYB_48__5_,
         u5_mult_82_CARRYB_48__6_, u5_mult_82_CARRYB_48__7_,
         u5_mult_82_CARRYB_48__8_, u5_mult_82_CARRYB_48__9_,
         u5_mult_82_CARRYB_48__10_, u5_mult_82_CARRYB_48__11_,
         u5_mult_82_CARRYB_48__12_, u5_mult_82_CARRYB_48__13_,
         u5_mult_82_CARRYB_48__14_, u5_mult_82_CARRYB_48__15_,
         u5_mult_82_CARRYB_48__16_, u5_mult_82_CARRYB_48__17_,
         u5_mult_82_CARRYB_48__18_, u5_mult_82_CARRYB_48__19_,
         u5_mult_82_CARRYB_48__20_, u5_mult_82_CARRYB_48__21_,
         u5_mult_82_CARRYB_48__22_, u5_mult_82_CARRYB_48__23_,
         u5_mult_82_CARRYB_48__24_, u5_mult_82_CARRYB_48__25_,
         u5_mult_82_CARRYB_48__26_, u5_mult_82_CARRYB_48__27_,
         u5_mult_82_CARRYB_48__28_, u5_mult_82_CARRYB_48__29_,
         u5_mult_82_CARRYB_48__30_, u5_mult_82_CARRYB_48__31_,
         u5_mult_82_CARRYB_48__32_, u5_mult_82_CARRYB_48__33_,
         u5_mult_82_CARRYB_48__34_, u5_mult_82_CARRYB_48__35_,
         u5_mult_82_CARRYB_48__36_, u5_mult_82_CARRYB_48__37_,
         u5_mult_82_CARRYB_48__38_, u5_mult_82_CARRYB_48__39_,
         u5_mult_82_CARRYB_48__40_, u5_mult_82_CARRYB_48__41_,
         u5_mult_82_CARRYB_48__42_, u5_mult_82_CARRYB_48__43_,
         u5_mult_82_CARRYB_48__44_, u5_mult_82_CARRYB_48__45_,
         u5_mult_82_CARRYB_48__46_, u5_mult_82_CARRYB_48__47_,
         u5_mult_82_CARRYB_48__48_, u5_mult_82_CARRYB_48__49_,
         u5_mult_82_CARRYB_48__50_, u5_mult_82_CARRYB_48__51_,
         u5_mult_82_CARRYB_49__0_, u5_mult_82_CARRYB_49__1_,
         u5_mult_82_CARRYB_49__2_, u5_mult_82_CARRYB_49__3_,
         u5_mult_82_CARRYB_49__4_, u5_mult_82_CARRYB_49__5_,
         u5_mult_82_CARRYB_49__6_, u5_mult_82_CARRYB_49__7_,
         u5_mult_82_CARRYB_49__8_, u5_mult_82_CARRYB_49__9_,
         u5_mult_82_CARRYB_49__10_, u5_mult_82_CARRYB_49__11_,
         u5_mult_82_CARRYB_49__12_, u5_mult_82_CARRYB_49__13_,
         u5_mult_82_CARRYB_49__14_, u5_mult_82_CARRYB_49__15_,
         u5_mult_82_CARRYB_49__16_, u5_mult_82_CARRYB_49__17_,
         u5_mult_82_CARRYB_49__18_, u5_mult_82_CARRYB_49__19_,
         u5_mult_82_CARRYB_49__20_, u5_mult_82_CARRYB_49__21_,
         u5_mult_82_CARRYB_49__22_, u5_mult_82_CARRYB_49__23_,
         u5_mult_82_CARRYB_49__24_, u5_mult_82_CARRYB_49__25_,
         u5_mult_82_CARRYB_49__26_, u5_mult_82_CARRYB_49__27_,
         u5_mult_82_CARRYB_49__28_, u5_mult_82_CARRYB_49__29_,
         u5_mult_82_CARRYB_49__30_, u5_mult_82_CARRYB_49__31_,
         u5_mult_82_CARRYB_49__32_, u5_mult_82_CARRYB_49__33_,
         u5_mult_82_CARRYB_49__34_, u5_mult_82_CARRYB_49__35_,
         u5_mult_82_CARRYB_49__36_, u5_mult_82_CARRYB_49__37_,
         u5_mult_82_CARRYB_49__38_, u5_mult_82_CARRYB_49__39_,
         u5_mult_82_CARRYB_49__40_, u5_mult_82_CARRYB_49__41_,
         u5_mult_82_CARRYB_49__42_, u5_mult_82_CARRYB_49__43_,
         u5_mult_82_CARRYB_49__44_, u5_mult_82_CARRYB_49__45_,
         u5_mult_82_CARRYB_49__46_, u5_mult_82_CARRYB_49__47_,
         u5_mult_82_CARRYB_49__48_, u5_mult_82_CARRYB_49__49_,
         u5_mult_82_CARRYB_49__50_, u5_mult_82_CARRYB_49__51_,
         u5_mult_82_CARRYB_50__0_, u5_mult_82_CARRYB_50__1_,
         u5_mult_82_CARRYB_50__2_, u5_mult_82_CARRYB_50__3_,
         u5_mult_82_CARRYB_50__4_, u5_mult_82_CARRYB_50__5_,
         u5_mult_82_CARRYB_50__6_, u5_mult_82_CARRYB_50__7_,
         u5_mult_82_CARRYB_50__8_, u5_mult_82_CARRYB_50__9_,
         u5_mult_82_CARRYB_50__10_, u5_mult_82_CARRYB_50__11_,
         u5_mult_82_CARRYB_50__12_, u5_mult_82_CARRYB_50__13_,
         u5_mult_82_CARRYB_50__14_, u5_mult_82_CARRYB_50__15_,
         u5_mult_82_CARRYB_50__16_, u5_mult_82_CARRYB_50__17_,
         u5_mult_82_CARRYB_50__18_, u5_mult_82_CARRYB_50__19_,
         u5_mult_82_CARRYB_50__20_, u5_mult_82_CARRYB_50__21_,
         u5_mult_82_CARRYB_50__22_, u5_mult_82_CARRYB_50__23_,
         u5_mult_82_CARRYB_50__24_, u5_mult_82_CARRYB_50__25_,
         u5_mult_82_CARRYB_50__26_, u5_mult_82_CARRYB_50__27_,
         u5_mult_82_CARRYB_50__28_, u5_mult_82_CARRYB_50__29_,
         u5_mult_82_CARRYB_50__30_, u5_mult_82_CARRYB_50__31_,
         u5_mult_82_CARRYB_50__32_, u5_mult_82_CARRYB_50__33_,
         u5_mult_82_CARRYB_50__34_, u5_mult_82_CARRYB_50__35_,
         u5_mult_82_CARRYB_50__36_, u5_mult_82_CARRYB_50__37_,
         u5_mult_82_CARRYB_50__38_, u5_mult_82_CARRYB_50__39_,
         u5_mult_82_CARRYB_50__40_, u5_mult_82_CARRYB_50__41_,
         u5_mult_82_CARRYB_50__42_, u5_mult_82_CARRYB_50__43_,
         u5_mult_82_CARRYB_50__44_, u5_mult_82_CARRYB_50__45_,
         u5_mult_82_CARRYB_50__46_, u5_mult_82_CARRYB_50__47_,
         u5_mult_82_CARRYB_50__48_, u5_mult_82_CARRYB_50__49_,
         u5_mult_82_CARRYB_50__50_, u5_mult_82_CARRYB_50__51_,
         u5_mult_82_CARRYB_51__0_, u5_mult_82_CARRYB_51__1_,
         u5_mult_82_CARRYB_51__2_, u5_mult_82_CARRYB_51__3_,
         u5_mult_82_CARRYB_51__4_, u5_mult_82_CARRYB_51__5_,
         u5_mult_82_CARRYB_51__6_, u5_mult_82_CARRYB_51__7_,
         u5_mult_82_CARRYB_51__8_, u5_mult_82_CARRYB_51__9_,
         u5_mult_82_CARRYB_51__10_, u5_mult_82_CARRYB_51__11_,
         u5_mult_82_CARRYB_51__12_, u5_mult_82_CARRYB_51__13_,
         u5_mult_82_CARRYB_51__14_, u5_mult_82_CARRYB_51__15_,
         u5_mult_82_CARRYB_51__16_, u5_mult_82_CARRYB_51__17_,
         u5_mult_82_CARRYB_51__18_, u5_mult_82_CARRYB_51__19_,
         u5_mult_82_CARRYB_51__20_, u5_mult_82_CARRYB_51__21_,
         u5_mult_82_CARRYB_51__22_, u5_mult_82_CARRYB_51__23_,
         u5_mult_82_CARRYB_51__24_, u5_mult_82_CARRYB_51__25_,
         u5_mult_82_CARRYB_51__26_, u5_mult_82_CARRYB_51__27_,
         u5_mult_82_CARRYB_51__28_, u5_mult_82_CARRYB_51__29_,
         u5_mult_82_CARRYB_51__30_, u5_mult_82_CARRYB_51__31_,
         u5_mult_82_CARRYB_51__32_, u5_mult_82_CARRYB_51__33_,
         u5_mult_82_CARRYB_51__34_, u5_mult_82_CARRYB_51__35_,
         u5_mult_82_CARRYB_51__36_, u5_mult_82_CARRYB_51__37_,
         u5_mult_82_CARRYB_51__38_, u5_mult_82_CARRYB_51__39_,
         u5_mult_82_CARRYB_51__40_, u5_mult_82_CARRYB_51__41_,
         u5_mult_82_CARRYB_51__42_, u5_mult_82_CARRYB_51__43_,
         u5_mult_82_CARRYB_51__44_, u5_mult_82_CARRYB_51__45_,
         u5_mult_82_CARRYB_51__46_, u5_mult_82_CARRYB_51__47_,
         u5_mult_82_CARRYB_51__48_, u5_mult_82_CARRYB_51__49_,
         u5_mult_82_CARRYB_51__50_, u5_mult_82_CARRYB_51__51_,
         u5_mult_82_CARRYB_52__0_, u5_mult_82_CARRYB_52__1_,
         u5_mult_82_CARRYB_52__2_, u5_mult_82_CARRYB_52__3_,
         u5_mult_82_CARRYB_52__4_, u5_mult_82_CARRYB_52__5_,
         u5_mult_82_CARRYB_52__6_, u5_mult_82_CARRYB_52__7_,
         u5_mult_82_CARRYB_52__8_, u5_mult_82_CARRYB_52__9_,
         u5_mult_82_CARRYB_52__10_, u5_mult_82_CARRYB_52__11_,
         u5_mult_82_CARRYB_52__12_, u5_mult_82_CARRYB_52__13_,
         u5_mult_82_CARRYB_52__14_, u5_mult_82_CARRYB_52__15_,
         u5_mult_82_CARRYB_52__16_, u5_mult_82_CARRYB_52__17_,
         u5_mult_82_CARRYB_52__18_, u5_mult_82_CARRYB_52__19_,
         u5_mult_82_CARRYB_52__20_, u5_mult_82_CARRYB_52__21_,
         u5_mult_82_CARRYB_52__22_, u5_mult_82_CARRYB_52__23_,
         u5_mult_82_CARRYB_52__24_, u5_mult_82_CARRYB_52__25_,
         u5_mult_82_CARRYB_52__26_, u5_mult_82_CARRYB_52__27_,
         u5_mult_82_CARRYB_52__28_, u5_mult_82_CARRYB_52__29_,
         u5_mult_82_CARRYB_52__30_, u5_mult_82_CARRYB_52__31_,
         u5_mult_82_CARRYB_52__32_, u5_mult_82_CARRYB_52__33_,
         u5_mult_82_CARRYB_52__34_, u5_mult_82_CARRYB_52__35_,
         u5_mult_82_CARRYB_52__36_, u5_mult_82_CARRYB_52__37_,
         u5_mult_82_CARRYB_52__38_, u5_mult_82_CARRYB_52__39_,
         u5_mult_82_CARRYB_52__40_, u5_mult_82_CARRYB_52__41_,
         u5_mult_82_CARRYB_52__42_, u5_mult_82_CARRYB_52__43_,
         u5_mult_82_CARRYB_52__44_, u5_mult_82_CARRYB_52__45_,
         u5_mult_82_CARRYB_52__46_, u5_mult_82_CARRYB_52__47_,
         u5_mult_82_CARRYB_52__48_, u5_mult_82_CARRYB_52__49_,
         u5_mult_82_CARRYB_52__50_, u5_mult_82_CARRYB_52__51_,
         u5_mult_82_SUMB_33__36_, u5_mult_82_SUMB_33__37_,
         u5_mult_82_SUMB_33__38_, u5_mult_82_SUMB_33__39_,
         u5_mult_82_SUMB_33__40_, u5_mult_82_SUMB_33__41_,
         u5_mult_82_SUMB_33__42_, u5_mult_82_SUMB_33__43_,
         u5_mult_82_SUMB_33__44_, u5_mult_82_SUMB_33__45_,
         u5_mult_82_SUMB_33__46_, u5_mult_82_SUMB_33__47_,
         u5_mult_82_SUMB_33__48_, u5_mult_82_SUMB_33__49_,
         u5_mult_82_SUMB_33__50_, u5_mult_82_SUMB_33__51_,
         u5_mult_82_SUMB_34__1_, u5_mult_82_SUMB_34__2_,
         u5_mult_82_SUMB_34__3_, u5_mult_82_SUMB_34__4_,
         u5_mult_82_SUMB_34__5_, u5_mult_82_SUMB_34__6_,
         u5_mult_82_SUMB_34__7_, u5_mult_82_SUMB_34__8_,
         u5_mult_82_SUMB_34__9_, u5_mult_82_SUMB_34__10_,
         u5_mult_82_SUMB_34__11_, u5_mult_82_SUMB_34__12_,
         u5_mult_82_SUMB_34__13_, u5_mult_82_SUMB_34__14_,
         u5_mult_82_SUMB_34__15_, u5_mult_82_SUMB_34__16_,
         u5_mult_82_SUMB_34__17_, u5_mult_82_SUMB_34__18_,
         u5_mult_82_SUMB_34__19_, u5_mult_82_SUMB_34__20_,
         u5_mult_82_SUMB_34__21_, u5_mult_82_SUMB_34__22_,
         u5_mult_82_SUMB_34__23_, u5_mult_82_SUMB_34__24_,
         u5_mult_82_SUMB_34__25_, u5_mult_82_SUMB_34__26_,
         u5_mult_82_SUMB_34__27_, u5_mult_82_SUMB_34__28_,
         u5_mult_82_SUMB_34__29_, u5_mult_82_SUMB_34__30_,
         u5_mult_82_SUMB_34__31_, u5_mult_82_SUMB_34__32_,
         u5_mult_82_SUMB_34__33_, u5_mult_82_SUMB_34__34_,
         u5_mult_82_SUMB_34__35_, u5_mult_82_SUMB_34__36_,
         u5_mult_82_SUMB_34__37_, u5_mult_82_SUMB_34__38_,
         u5_mult_82_SUMB_34__39_, u5_mult_82_SUMB_34__40_,
         u5_mult_82_SUMB_34__41_, u5_mult_82_SUMB_34__42_,
         u5_mult_82_SUMB_34__43_, u5_mult_82_SUMB_34__44_,
         u5_mult_82_SUMB_34__45_, u5_mult_82_SUMB_34__46_,
         u5_mult_82_SUMB_34__47_, u5_mult_82_SUMB_34__48_,
         u5_mult_82_SUMB_34__49_, u5_mult_82_SUMB_34__50_,
         u5_mult_82_SUMB_34__51_, u5_mult_82_SUMB_35__1_,
         u5_mult_82_SUMB_35__2_, u5_mult_82_SUMB_35__3_,
         u5_mult_82_SUMB_35__4_, u5_mult_82_SUMB_35__5_,
         u5_mult_82_SUMB_35__6_, u5_mult_82_SUMB_35__7_,
         u5_mult_82_SUMB_35__8_, u5_mult_82_SUMB_35__9_,
         u5_mult_82_SUMB_35__10_, u5_mult_82_SUMB_35__11_,
         u5_mult_82_SUMB_35__12_, u5_mult_82_SUMB_35__13_,
         u5_mult_82_SUMB_35__14_, u5_mult_82_SUMB_35__15_,
         u5_mult_82_SUMB_35__16_, u5_mult_82_SUMB_35__17_,
         u5_mult_82_SUMB_35__18_, u5_mult_82_SUMB_35__19_,
         u5_mult_82_SUMB_35__20_, u5_mult_82_SUMB_35__21_,
         u5_mult_82_SUMB_35__22_, u5_mult_82_SUMB_35__23_,
         u5_mult_82_SUMB_35__24_, u5_mult_82_SUMB_35__25_,
         u5_mult_82_SUMB_35__26_, u5_mult_82_SUMB_35__27_,
         u5_mult_82_SUMB_35__28_, u5_mult_82_SUMB_35__29_,
         u5_mult_82_SUMB_35__30_, u5_mult_82_SUMB_35__31_,
         u5_mult_82_SUMB_35__32_, u5_mult_82_SUMB_35__33_,
         u5_mult_82_SUMB_35__34_, u5_mult_82_SUMB_35__35_,
         u5_mult_82_SUMB_35__36_, u5_mult_82_SUMB_35__37_,
         u5_mult_82_SUMB_35__38_, u5_mult_82_SUMB_35__39_,
         u5_mult_82_SUMB_35__40_, u5_mult_82_SUMB_35__41_,
         u5_mult_82_SUMB_35__42_, u5_mult_82_SUMB_35__43_,
         u5_mult_82_SUMB_35__44_, u5_mult_82_SUMB_35__45_,
         u5_mult_82_SUMB_35__46_, u5_mult_82_SUMB_35__47_,
         u5_mult_82_SUMB_35__48_, u5_mult_82_SUMB_35__49_,
         u5_mult_82_SUMB_35__50_, u5_mult_82_SUMB_35__51_,
         u5_mult_82_SUMB_36__1_, u5_mult_82_SUMB_36__2_,
         u5_mult_82_SUMB_36__3_, u5_mult_82_SUMB_36__4_,
         u5_mult_82_SUMB_36__5_, u5_mult_82_SUMB_36__6_,
         u5_mult_82_SUMB_36__7_, u5_mult_82_SUMB_36__8_,
         u5_mult_82_SUMB_36__9_, u5_mult_82_SUMB_36__10_,
         u5_mult_82_SUMB_36__11_, u5_mult_82_SUMB_36__12_,
         u5_mult_82_SUMB_36__13_, u5_mult_82_SUMB_36__14_,
         u5_mult_82_SUMB_36__15_, u5_mult_82_SUMB_36__16_,
         u5_mult_82_SUMB_36__17_, u5_mult_82_SUMB_36__18_,
         u5_mult_82_SUMB_36__19_, u5_mult_82_SUMB_36__20_,
         u5_mult_82_SUMB_36__21_, u5_mult_82_SUMB_36__22_,
         u5_mult_82_SUMB_36__23_, u5_mult_82_SUMB_36__24_,
         u5_mult_82_SUMB_36__25_, u5_mult_82_SUMB_36__26_,
         u5_mult_82_SUMB_36__27_, u5_mult_82_SUMB_36__28_,
         u5_mult_82_SUMB_36__29_, u5_mult_82_SUMB_36__30_,
         u5_mult_82_SUMB_36__31_, u5_mult_82_SUMB_36__32_,
         u5_mult_82_SUMB_36__33_, u5_mult_82_SUMB_36__34_,
         u5_mult_82_SUMB_36__35_, u5_mult_82_SUMB_36__36_,
         u5_mult_82_SUMB_36__37_, u5_mult_82_SUMB_36__38_,
         u5_mult_82_SUMB_36__39_, u5_mult_82_SUMB_36__40_,
         u5_mult_82_SUMB_36__41_, u5_mult_82_SUMB_36__42_,
         u5_mult_82_SUMB_36__43_, u5_mult_82_SUMB_36__44_,
         u5_mult_82_SUMB_36__45_, u5_mult_82_SUMB_36__46_,
         u5_mult_82_SUMB_36__47_, u5_mult_82_SUMB_36__48_,
         u5_mult_82_SUMB_36__49_, u5_mult_82_SUMB_36__50_,
         u5_mult_82_SUMB_36__51_, u5_mult_82_SUMB_37__1_,
         u5_mult_82_SUMB_37__2_, u5_mult_82_SUMB_37__3_,
         u5_mult_82_SUMB_37__4_, u5_mult_82_SUMB_37__5_,
         u5_mult_82_SUMB_37__6_, u5_mult_82_SUMB_37__7_,
         u5_mult_82_SUMB_37__8_, u5_mult_82_SUMB_37__9_,
         u5_mult_82_SUMB_37__10_, u5_mult_82_SUMB_37__11_,
         u5_mult_82_SUMB_37__12_, u5_mult_82_SUMB_37__13_,
         u5_mult_82_SUMB_37__14_, u5_mult_82_SUMB_37__15_,
         u5_mult_82_SUMB_37__16_, u5_mult_82_SUMB_37__17_,
         u5_mult_82_SUMB_37__18_, u5_mult_82_SUMB_37__19_,
         u5_mult_82_SUMB_37__20_, u5_mult_82_SUMB_37__21_,
         u5_mult_82_SUMB_37__22_, u5_mult_82_SUMB_37__23_,
         u5_mult_82_SUMB_37__24_, u5_mult_82_SUMB_37__25_,
         u5_mult_82_SUMB_37__26_, u5_mult_82_SUMB_37__27_,
         u5_mult_82_SUMB_37__28_, u5_mult_82_SUMB_37__29_,
         u5_mult_82_SUMB_37__30_, u5_mult_82_SUMB_37__31_,
         u5_mult_82_SUMB_37__32_, u5_mult_82_SUMB_37__33_,
         u5_mult_82_SUMB_37__34_, u5_mult_82_SUMB_37__35_,
         u5_mult_82_SUMB_37__36_, u5_mult_82_SUMB_37__37_,
         u5_mult_82_SUMB_37__38_, u5_mult_82_SUMB_37__39_,
         u5_mult_82_SUMB_37__40_, u5_mult_82_SUMB_37__41_,
         u5_mult_82_SUMB_37__42_, u5_mult_82_SUMB_37__43_,
         u5_mult_82_SUMB_37__44_, u5_mult_82_SUMB_37__45_,
         u5_mult_82_SUMB_37__46_, u5_mult_82_SUMB_37__47_,
         u5_mult_82_SUMB_37__48_, u5_mult_82_SUMB_37__49_,
         u5_mult_82_SUMB_37__50_, u5_mult_82_SUMB_37__51_,
         u5_mult_82_SUMB_38__1_, u5_mult_82_SUMB_38__2_,
         u5_mult_82_SUMB_38__3_, u5_mult_82_SUMB_38__4_,
         u5_mult_82_SUMB_38__5_, u5_mult_82_SUMB_38__6_,
         u5_mult_82_SUMB_38__7_, u5_mult_82_SUMB_38__8_,
         u5_mult_82_SUMB_38__9_, u5_mult_82_SUMB_38__10_,
         u5_mult_82_SUMB_38__11_, u5_mult_82_SUMB_38__12_,
         u5_mult_82_SUMB_38__13_, u5_mult_82_SUMB_38__14_,
         u5_mult_82_SUMB_38__15_, u5_mult_82_SUMB_38__16_,
         u5_mult_82_SUMB_38__17_, u5_mult_82_SUMB_38__18_,
         u5_mult_82_SUMB_38__19_, u5_mult_82_SUMB_38__20_,
         u5_mult_82_SUMB_38__21_, u5_mult_82_SUMB_38__22_,
         u5_mult_82_SUMB_38__23_, u5_mult_82_SUMB_38__24_,
         u5_mult_82_SUMB_38__25_, u5_mult_82_SUMB_38__26_,
         u5_mult_82_SUMB_38__27_, u5_mult_82_SUMB_38__28_,
         u5_mult_82_SUMB_38__29_, u5_mult_82_SUMB_38__30_,
         u5_mult_82_SUMB_38__31_, u5_mult_82_SUMB_38__32_,
         u5_mult_82_SUMB_38__33_, u5_mult_82_SUMB_38__34_,
         u5_mult_82_SUMB_38__35_, u5_mult_82_SUMB_38__36_,
         u5_mult_82_SUMB_38__37_, u5_mult_82_SUMB_38__38_,
         u5_mult_82_SUMB_38__39_, u5_mult_82_SUMB_38__40_,
         u5_mult_82_SUMB_38__41_, u5_mult_82_SUMB_38__42_,
         u5_mult_82_SUMB_38__43_, u5_mult_82_SUMB_38__44_,
         u5_mult_82_SUMB_38__45_, u5_mult_82_SUMB_38__46_,
         u5_mult_82_SUMB_38__47_, u5_mult_82_SUMB_38__48_,
         u5_mult_82_SUMB_38__49_, u5_mult_82_SUMB_38__50_,
         u5_mult_82_SUMB_38__51_, u5_mult_82_SUMB_39__1_,
         u5_mult_82_SUMB_39__2_, u5_mult_82_SUMB_39__3_,
         u5_mult_82_SUMB_39__4_, u5_mult_82_SUMB_39__5_,
         u5_mult_82_SUMB_39__6_, u5_mult_82_SUMB_39__7_,
         u5_mult_82_SUMB_39__8_, u5_mult_82_SUMB_39__9_,
         u5_mult_82_SUMB_39__10_, u5_mult_82_SUMB_39__11_,
         u5_mult_82_SUMB_39__12_, u5_mult_82_SUMB_39__13_,
         u5_mult_82_SUMB_39__14_, u5_mult_82_SUMB_39__15_,
         u5_mult_82_SUMB_39__16_, u5_mult_82_SUMB_39__17_,
         u5_mult_82_SUMB_39__18_, u5_mult_82_SUMB_39__19_,
         u5_mult_82_SUMB_39__20_, u5_mult_82_SUMB_39__21_,
         u5_mult_82_SUMB_39__22_, u5_mult_82_SUMB_39__23_,
         u5_mult_82_SUMB_39__24_, u5_mult_82_SUMB_39__25_,
         u5_mult_82_SUMB_39__26_, u5_mult_82_SUMB_39__27_,
         u5_mult_82_SUMB_39__28_, u5_mult_82_SUMB_39__29_,
         u5_mult_82_SUMB_39__30_, u5_mult_82_SUMB_39__31_,
         u5_mult_82_SUMB_39__32_, u5_mult_82_SUMB_39__33_,
         u5_mult_82_SUMB_39__34_, u5_mult_82_SUMB_39__35_,
         u5_mult_82_SUMB_39__36_, u5_mult_82_SUMB_39__37_,
         u5_mult_82_SUMB_39__38_, u5_mult_82_SUMB_39__39_,
         u5_mult_82_SUMB_39__40_, u5_mult_82_SUMB_39__41_,
         u5_mult_82_SUMB_39__42_, u5_mult_82_SUMB_39__43_,
         u5_mult_82_SUMB_39__44_, u5_mult_82_SUMB_39__45_,
         u5_mult_82_SUMB_39__46_, u5_mult_82_SUMB_39__47_,
         u5_mult_82_SUMB_39__48_, u5_mult_82_SUMB_39__49_,
         u5_mult_82_SUMB_39__50_, u5_mult_82_SUMB_39__51_,
         u5_mult_82_SUMB_40__1_, u5_mult_82_SUMB_40__2_,
         u5_mult_82_SUMB_40__3_, u5_mult_82_SUMB_40__4_,
         u5_mult_82_SUMB_40__5_, u5_mult_82_SUMB_40__6_,
         u5_mult_82_SUMB_40__7_, u5_mult_82_SUMB_40__8_,
         u5_mult_82_SUMB_40__9_, u5_mult_82_SUMB_40__10_,
         u5_mult_82_SUMB_40__11_, u5_mult_82_SUMB_40__12_,
         u5_mult_82_SUMB_40__13_, u5_mult_82_SUMB_40__14_,
         u5_mult_82_SUMB_40__15_, u5_mult_82_SUMB_40__16_,
         u5_mult_82_SUMB_40__17_, u5_mult_82_SUMB_40__18_,
         u5_mult_82_SUMB_40__19_, u5_mult_82_SUMB_40__20_,
         u5_mult_82_SUMB_40__21_, u5_mult_82_SUMB_40__22_,
         u5_mult_82_SUMB_40__23_, u5_mult_82_SUMB_40__24_,
         u5_mult_82_SUMB_40__25_, u5_mult_82_SUMB_40__26_,
         u5_mult_82_SUMB_40__27_, u5_mult_82_SUMB_40__28_,
         u5_mult_82_SUMB_40__29_, u5_mult_82_SUMB_40__30_,
         u5_mult_82_SUMB_40__31_, u5_mult_82_SUMB_40__32_,
         u5_mult_82_SUMB_40__33_, u5_mult_82_SUMB_40__34_,
         u5_mult_82_SUMB_40__35_, u5_mult_82_SUMB_40__36_,
         u5_mult_82_SUMB_40__37_, u5_mult_82_SUMB_40__38_,
         u5_mult_82_SUMB_40__39_, u5_mult_82_SUMB_40__40_,
         u5_mult_82_SUMB_40__41_, u5_mult_82_SUMB_40__42_,
         u5_mult_82_SUMB_40__43_, u5_mult_82_SUMB_40__44_,
         u5_mult_82_SUMB_40__45_, u5_mult_82_SUMB_40__46_,
         u5_mult_82_SUMB_40__47_, u5_mult_82_SUMB_40__48_,
         u5_mult_82_SUMB_40__49_, u5_mult_82_SUMB_40__50_,
         u5_mult_82_SUMB_40__51_, u5_mult_82_SUMB_41__1_,
         u5_mult_82_SUMB_41__2_, u5_mult_82_SUMB_41__3_,
         u5_mult_82_SUMB_41__4_, u5_mult_82_SUMB_41__5_,
         u5_mult_82_SUMB_41__6_, u5_mult_82_SUMB_41__7_,
         u5_mult_82_SUMB_41__8_, u5_mult_82_SUMB_41__9_,
         u5_mult_82_SUMB_41__10_, u5_mult_82_SUMB_41__11_,
         u5_mult_82_SUMB_41__12_, u5_mult_82_SUMB_41__13_,
         u5_mult_82_SUMB_41__14_, u5_mult_82_SUMB_41__15_,
         u5_mult_82_SUMB_41__16_, u5_mult_82_SUMB_41__17_,
         u5_mult_82_SUMB_41__18_, u5_mult_82_SUMB_41__19_,
         u5_mult_82_SUMB_41__20_, u5_mult_82_SUMB_41__21_,
         u5_mult_82_SUMB_41__22_, u5_mult_82_SUMB_41__23_,
         u5_mult_82_SUMB_41__24_, u5_mult_82_SUMB_41__25_,
         u5_mult_82_SUMB_41__26_, u5_mult_82_SUMB_41__27_,
         u5_mult_82_SUMB_41__28_, u5_mult_82_SUMB_41__29_,
         u5_mult_82_SUMB_41__30_, u5_mult_82_SUMB_41__31_,
         u5_mult_82_SUMB_41__32_, u5_mult_82_SUMB_41__33_,
         u5_mult_82_SUMB_41__34_, u5_mult_82_SUMB_41__35_,
         u5_mult_82_SUMB_41__36_, u5_mult_82_SUMB_41__37_,
         u5_mult_82_SUMB_41__38_, u5_mult_82_SUMB_41__39_,
         u5_mult_82_SUMB_41__40_, u5_mult_82_SUMB_41__41_,
         u5_mult_82_SUMB_41__42_, u5_mult_82_SUMB_41__43_,
         u5_mult_82_SUMB_41__44_, u5_mult_82_SUMB_41__45_,
         u5_mult_82_SUMB_41__46_, u5_mult_82_SUMB_41__47_,
         u5_mult_82_SUMB_41__48_, u5_mult_82_SUMB_41__49_,
         u5_mult_82_SUMB_41__50_, u5_mult_82_SUMB_41__51_,
         u5_mult_82_SUMB_42__1_, u5_mult_82_SUMB_42__2_,
         u5_mult_82_SUMB_42__3_, u5_mult_82_SUMB_42__4_,
         u5_mult_82_SUMB_42__5_, u5_mult_82_SUMB_42__6_,
         u5_mult_82_SUMB_42__7_, u5_mult_82_SUMB_42__8_,
         u5_mult_82_SUMB_42__9_, u5_mult_82_SUMB_42__10_,
         u5_mult_82_SUMB_42__11_, u5_mult_82_SUMB_42__12_,
         u5_mult_82_SUMB_42__13_, u5_mult_82_SUMB_42__14_,
         u5_mult_82_SUMB_42__15_, u5_mult_82_SUMB_42__16_,
         u5_mult_82_SUMB_42__17_, u5_mult_82_SUMB_42__18_,
         u5_mult_82_SUMB_42__19_, u5_mult_82_SUMB_42__20_,
         u5_mult_82_SUMB_42__21_, u5_mult_82_SUMB_42__22_,
         u5_mult_82_SUMB_42__23_, u5_mult_82_SUMB_42__24_,
         u5_mult_82_SUMB_42__25_, u5_mult_82_SUMB_42__26_,
         u5_mult_82_SUMB_42__27_, u5_mult_82_SUMB_42__28_,
         u5_mult_82_SUMB_42__29_, u5_mult_82_SUMB_42__30_,
         u5_mult_82_SUMB_42__31_, u5_mult_82_SUMB_42__32_,
         u5_mult_82_SUMB_42__33_, u5_mult_82_SUMB_42__34_,
         u5_mult_82_SUMB_42__35_, u5_mult_82_SUMB_42__36_,
         u5_mult_82_SUMB_42__37_, u5_mult_82_SUMB_42__38_,
         u5_mult_82_SUMB_42__39_, u5_mult_82_SUMB_42__40_,
         u5_mult_82_SUMB_42__41_, u5_mult_82_SUMB_42__42_,
         u5_mult_82_SUMB_42__43_, u5_mult_82_SUMB_42__44_,
         u5_mult_82_SUMB_42__45_, u5_mult_82_SUMB_42__46_,
         u5_mult_82_SUMB_42__47_, u5_mult_82_SUMB_42__48_,
         u5_mult_82_SUMB_42__49_, u5_mult_82_SUMB_42__50_,
         u5_mult_82_SUMB_42__51_, u5_mult_82_SUMB_43__1_,
         u5_mult_82_SUMB_43__2_, u5_mult_82_SUMB_43__3_,
         u5_mult_82_SUMB_43__4_, u5_mult_82_SUMB_43__5_,
         u5_mult_82_SUMB_43__6_, u5_mult_82_SUMB_43__7_,
         u5_mult_82_SUMB_43__8_, u5_mult_82_SUMB_43__9_,
         u5_mult_82_SUMB_43__10_, u5_mult_82_SUMB_43__11_,
         u5_mult_82_SUMB_43__12_, u5_mult_82_SUMB_43__13_,
         u5_mult_82_SUMB_43__14_, u5_mult_82_SUMB_43__15_,
         u5_mult_82_SUMB_43__16_, u5_mult_82_SUMB_43__17_,
         u5_mult_82_CARRYB_33__36_, u5_mult_82_CARRYB_33__37_,
         u5_mult_82_CARRYB_33__38_, u5_mult_82_CARRYB_33__39_,
         u5_mult_82_CARRYB_33__40_, u5_mult_82_CARRYB_33__41_,
         u5_mult_82_CARRYB_33__42_, u5_mult_82_CARRYB_33__43_,
         u5_mult_82_CARRYB_33__44_, u5_mult_82_CARRYB_33__45_,
         u5_mult_82_CARRYB_33__46_, u5_mult_82_CARRYB_33__47_,
         u5_mult_82_CARRYB_33__48_, u5_mult_82_CARRYB_33__49_,
         u5_mult_82_CARRYB_33__50_, u5_mult_82_CARRYB_33__51_,
         u5_mult_82_CARRYB_34__0_, u5_mult_82_CARRYB_34__1_,
         u5_mult_82_CARRYB_34__2_, u5_mult_82_CARRYB_34__3_,
         u5_mult_82_CARRYB_34__4_, u5_mult_82_CARRYB_34__5_,
         u5_mult_82_CARRYB_34__6_, u5_mult_82_CARRYB_34__7_,
         u5_mult_82_CARRYB_34__8_, u5_mult_82_CARRYB_34__9_,
         u5_mult_82_CARRYB_34__10_, u5_mult_82_CARRYB_34__11_,
         u5_mult_82_CARRYB_34__12_, u5_mult_82_CARRYB_34__13_,
         u5_mult_82_CARRYB_34__14_, u5_mult_82_CARRYB_34__15_,
         u5_mult_82_CARRYB_34__16_, u5_mult_82_CARRYB_34__17_,
         u5_mult_82_CARRYB_34__18_, u5_mult_82_CARRYB_34__19_,
         u5_mult_82_CARRYB_34__20_, u5_mult_82_CARRYB_34__21_,
         u5_mult_82_CARRYB_34__22_, u5_mult_82_CARRYB_34__23_,
         u5_mult_82_CARRYB_34__24_, u5_mult_82_CARRYB_34__25_,
         u5_mult_82_CARRYB_34__26_, u5_mult_82_CARRYB_34__27_,
         u5_mult_82_CARRYB_34__28_, u5_mult_82_CARRYB_34__29_,
         u5_mult_82_CARRYB_34__30_, u5_mult_82_CARRYB_34__31_,
         u5_mult_82_CARRYB_34__32_, u5_mult_82_CARRYB_34__33_,
         u5_mult_82_CARRYB_34__34_, u5_mult_82_CARRYB_34__35_,
         u5_mult_82_CARRYB_34__36_, u5_mult_82_CARRYB_34__37_,
         u5_mult_82_CARRYB_34__38_, u5_mult_82_CARRYB_34__39_,
         u5_mult_82_CARRYB_34__40_, u5_mult_82_CARRYB_34__41_,
         u5_mult_82_CARRYB_34__42_, u5_mult_82_CARRYB_34__43_,
         u5_mult_82_CARRYB_34__44_, u5_mult_82_CARRYB_34__45_,
         u5_mult_82_CARRYB_34__46_, u5_mult_82_CARRYB_34__47_,
         u5_mult_82_CARRYB_34__48_, u5_mult_82_CARRYB_34__49_,
         u5_mult_82_CARRYB_34__50_, u5_mult_82_CARRYB_34__51_,
         u5_mult_82_CARRYB_35__0_, u5_mult_82_CARRYB_35__1_,
         u5_mult_82_CARRYB_35__2_, u5_mult_82_CARRYB_35__3_,
         u5_mult_82_CARRYB_35__4_, u5_mult_82_CARRYB_35__5_,
         u5_mult_82_CARRYB_35__6_, u5_mult_82_CARRYB_35__7_,
         u5_mult_82_CARRYB_35__8_, u5_mult_82_CARRYB_35__9_,
         u5_mult_82_CARRYB_35__10_, u5_mult_82_CARRYB_35__11_,
         u5_mult_82_CARRYB_35__12_, u5_mult_82_CARRYB_35__13_,
         u5_mult_82_CARRYB_35__14_, u5_mult_82_CARRYB_35__15_,
         u5_mult_82_CARRYB_35__16_, u5_mult_82_CARRYB_35__17_,
         u5_mult_82_CARRYB_35__18_, u5_mult_82_CARRYB_35__19_,
         u5_mult_82_CARRYB_35__20_, u5_mult_82_CARRYB_35__21_,
         u5_mult_82_CARRYB_35__22_, u5_mult_82_CARRYB_35__23_,
         u5_mult_82_CARRYB_35__24_, u5_mult_82_CARRYB_35__25_,
         u5_mult_82_CARRYB_35__26_, u5_mult_82_CARRYB_35__27_,
         u5_mult_82_CARRYB_35__28_, u5_mult_82_CARRYB_35__29_,
         u5_mult_82_CARRYB_35__30_, u5_mult_82_CARRYB_35__31_,
         u5_mult_82_CARRYB_35__32_, u5_mult_82_CARRYB_35__33_,
         u5_mult_82_CARRYB_35__34_, u5_mult_82_CARRYB_35__35_,
         u5_mult_82_CARRYB_35__36_, u5_mult_82_CARRYB_35__37_,
         u5_mult_82_CARRYB_35__38_, u5_mult_82_CARRYB_35__39_,
         u5_mult_82_CARRYB_35__40_, u5_mult_82_CARRYB_35__41_,
         u5_mult_82_CARRYB_35__42_, u5_mult_82_CARRYB_35__43_,
         u5_mult_82_CARRYB_35__44_, u5_mult_82_CARRYB_35__45_,
         u5_mult_82_CARRYB_35__46_, u5_mult_82_CARRYB_35__47_,
         u5_mult_82_CARRYB_35__48_, u5_mult_82_CARRYB_35__49_,
         u5_mult_82_CARRYB_35__50_, u5_mult_82_CARRYB_35__51_,
         u5_mult_82_CARRYB_36__0_, u5_mult_82_CARRYB_36__1_,
         u5_mult_82_CARRYB_36__2_, u5_mult_82_CARRYB_36__3_,
         u5_mult_82_CARRYB_36__4_, u5_mult_82_CARRYB_36__5_,
         u5_mult_82_CARRYB_36__6_, u5_mult_82_CARRYB_36__7_,
         u5_mult_82_CARRYB_36__8_, u5_mult_82_CARRYB_36__9_,
         u5_mult_82_CARRYB_36__10_, u5_mult_82_CARRYB_36__11_,
         u5_mult_82_CARRYB_36__12_, u5_mult_82_CARRYB_36__13_,
         u5_mult_82_CARRYB_36__14_, u5_mult_82_CARRYB_36__15_,
         u5_mult_82_CARRYB_36__16_, u5_mult_82_CARRYB_36__17_,
         u5_mult_82_CARRYB_36__18_, u5_mult_82_CARRYB_36__19_,
         u5_mult_82_CARRYB_36__20_, u5_mult_82_CARRYB_36__21_,
         u5_mult_82_CARRYB_36__22_, u5_mult_82_CARRYB_36__23_,
         u5_mult_82_CARRYB_36__24_, u5_mult_82_CARRYB_36__25_,
         u5_mult_82_CARRYB_36__26_, u5_mult_82_CARRYB_36__27_,
         u5_mult_82_CARRYB_36__28_, u5_mult_82_CARRYB_36__29_,
         u5_mult_82_CARRYB_36__30_, u5_mult_82_CARRYB_36__31_,
         u5_mult_82_CARRYB_36__32_, u5_mult_82_CARRYB_36__33_,
         u5_mult_82_CARRYB_36__34_, u5_mult_82_CARRYB_36__35_,
         u5_mult_82_CARRYB_36__36_, u5_mult_82_CARRYB_36__37_,
         u5_mult_82_CARRYB_36__38_, u5_mult_82_CARRYB_36__39_,
         u5_mult_82_CARRYB_36__40_, u5_mult_82_CARRYB_36__41_,
         u5_mult_82_CARRYB_36__42_, u5_mult_82_CARRYB_36__43_,
         u5_mult_82_CARRYB_36__44_, u5_mult_82_CARRYB_36__45_,
         u5_mult_82_CARRYB_36__46_, u5_mult_82_CARRYB_36__47_,
         u5_mult_82_CARRYB_36__48_, u5_mult_82_CARRYB_36__49_,
         u5_mult_82_CARRYB_36__50_, u5_mult_82_CARRYB_36__51_,
         u5_mult_82_CARRYB_37__0_, u5_mult_82_CARRYB_37__1_,
         u5_mult_82_CARRYB_37__2_, u5_mult_82_CARRYB_37__3_,
         u5_mult_82_CARRYB_37__4_, u5_mult_82_CARRYB_37__5_,
         u5_mult_82_CARRYB_37__6_, u5_mult_82_CARRYB_37__7_,
         u5_mult_82_CARRYB_37__8_, u5_mult_82_CARRYB_37__9_,
         u5_mult_82_CARRYB_37__10_, u5_mult_82_CARRYB_37__11_,
         u5_mult_82_CARRYB_37__12_, u5_mult_82_CARRYB_37__13_,
         u5_mult_82_CARRYB_37__14_, u5_mult_82_CARRYB_37__15_,
         u5_mult_82_CARRYB_37__16_, u5_mult_82_CARRYB_37__17_,
         u5_mult_82_CARRYB_37__18_, u5_mult_82_CARRYB_37__19_,
         u5_mult_82_CARRYB_37__20_, u5_mult_82_CARRYB_37__21_,
         u5_mult_82_CARRYB_37__22_, u5_mult_82_CARRYB_37__23_,
         u5_mult_82_CARRYB_37__24_, u5_mult_82_CARRYB_37__25_,
         u5_mult_82_CARRYB_37__26_, u5_mult_82_CARRYB_37__27_,
         u5_mult_82_CARRYB_37__28_, u5_mult_82_CARRYB_37__29_,
         u5_mult_82_CARRYB_37__30_, u5_mult_82_CARRYB_37__31_,
         u5_mult_82_CARRYB_37__32_, u5_mult_82_CARRYB_37__33_,
         u5_mult_82_CARRYB_37__34_, u5_mult_82_CARRYB_37__35_,
         u5_mult_82_CARRYB_37__36_, u5_mult_82_CARRYB_37__37_,
         u5_mult_82_CARRYB_37__38_, u5_mult_82_CARRYB_37__39_,
         u5_mult_82_CARRYB_37__40_, u5_mult_82_CARRYB_37__41_,
         u5_mult_82_CARRYB_37__42_, u5_mult_82_CARRYB_37__43_,
         u5_mult_82_CARRYB_37__44_, u5_mult_82_CARRYB_37__45_,
         u5_mult_82_CARRYB_37__46_, u5_mult_82_CARRYB_37__47_,
         u5_mult_82_CARRYB_37__48_, u5_mult_82_CARRYB_37__49_,
         u5_mult_82_CARRYB_37__50_, u5_mult_82_CARRYB_37__51_,
         u5_mult_82_CARRYB_38__0_, u5_mult_82_CARRYB_38__1_,
         u5_mult_82_CARRYB_38__2_, u5_mult_82_CARRYB_38__3_,
         u5_mult_82_CARRYB_38__4_, u5_mult_82_CARRYB_38__5_,
         u5_mult_82_CARRYB_38__6_, u5_mult_82_CARRYB_38__7_,
         u5_mult_82_CARRYB_38__8_, u5_mult_82_CARRYB_38__9_,
         u5_mult_82_CARRYB_38__10_, u5_mult_82_CARRYB_38__11_,
         u5_mult_82_CARRYB_38__12_, u5_mult_82_CARRYB_38__13_,
         u5_mult_82_CARRYB_38__14_, u5_mult_82_CARRYB_38__15_,
         u5_mult_82_CARRYB_38__16_, u5_mult_82_CARRYB_38__17_,
         u5_mult_82_CARRYB_38__18_, u5_mult_82_CARRYB_38__19_,
         u5_mult_82_CARRYB_38__20_, u5_mult_82_CARRYB_38__21_,
         u5_mult_82_CARRYB_38__22_, u5_mult_82_CARRYB_38__23_,
         u5_mult_82_CARRYB_38__24_, u5_mult_82_CARRYB_38__25_,
         u5_mult_82_CARRYB_38__26_, u5_mult_82_CARRYB_38__27_,
         u5_mult_82_CARRYB_38__28_, u5_mult_82_CARRYB_38__29_,
         u5_mult_82_CARRYB_38__30_, u5_mult_82_CARRYB_38__31_,
         u5_mult_82_CARRYB_38__32_, u5_mult_82_CARRYB_38__33_,
         u5_mult_82_CARRYB_38__34_, u5_mult_82_CARRYB_38__35_,
         u5_mult_82_CARRYB_38__36_, u5_mult_82_CARRYB_38__37_,
         u5_mult_82_CARRYB_38__38_, u5_mult_82_CARRYB_38__39_,
         u5_mult_82_CARRYB_38__40_, u5_mult_82_CARRYB_38__41_,
         u5_mult_82_CARRYB_38__42_, u5_mult_82_CARRYB_38__43_,
         u5_mult_82_CARRYB_38__44_, u5_mult_82_CARRYB_38__45_,
         u5_mult_82_CARRYB_38__46_, u5_mult_82_CARRYB_38__47_,
         u5_mult_82_CARRYB_38__48_, u5_mult_82_CARRYB_38__49_,
         u5_mult_82_CARRYB_38__50_, u5_mult_82_CARRYB_38__51_,
         u5_mult_82_CARRYB_39__0_, u5_mult_82_CARRYB_39__1_,
         u5_mult_82_CARRYB_39__2_, u5_mult_82_CARRYB_39__3_,
         u5_mult_82_CARRYB_39__4_, u5_mult_82_CARRYB_39__5_,
         u5_mult_82_CARRYB_39__6_, u5_mult_82_CARRYB_39__7_,
         u5_mult_82_CARRYB_39__8_, u5_mult_82_CARRYB_39__9_,
         u5_mult_82_CARRYB_39__10_, u5_mult_82_CARRYB_39__11_,
         u5_mult_82_CARRYB_39__12_, u5_mult_82_CARRYB_39__13_,
         u5_mult_82_CARRYB_39__14_, u5_mult_82_CARRYB_39__15_,
         u5_mult_82_CARRYB_39__16_, u5_mult_82_CARRYB_39__17_,
         u5_mult_82_CARRYB_39__18_, u5_mult_82_CARRYB_39__19_,
         u5_mult_82_CARRYB_39__20_, u5_mult_82_CARRYB_39__21_,
         u5_mult_82_CARRYB_39__22_, u5_mult_82_CARRYB_39__23_,
         u5_mult_82_CARRYB_39__24_, u5_mult_82_CARRYB_39__25_,
         u5_mult_82_CARRYB_39__26_, u5_mult_82_CARRYB_39__27_,
         u5_mult_82_CARRYB_39__28_, u5_mult_82_CARRYB_39__29_,
         u5_mult_82_CARRYB_39__30_, u5_mult_82_CARRYB_39__31_,
         u5_mult_82_CARRYB_39__32_, u5_mult_82_CARRYB_39__33_,
         u5_mult_82_CARRYB_39__34_, u5_mult_82_CARRYB_39__35_,
         u5_mult_82_CARRYB_39__36_, u5_mult_82_CARRYB_39__37_,
         u5_mult_82_CARRYB_39__38_, u5_mult_82_CARRYB_39__39_,
         u5_mult_82_CARRYB_39__40_, u5_mult_82_CARRYB_39__41_,
         u5_mult_82_CARRYB_39__42_, u5_mult_82_CARRYB_39__43_,
         u5_mult_82_CARRYB_39__44_, u5_mult_82_CARRYB_39__45_,
         u5_mult_82_CARRYB_39__46_, u5_mult_82_CARRYB_39__47_,
         u5_mult_82_CARRYB_39__48_, u5_mult_82_CARRYB_39__49_,
         u5_mult_82_CARRYB_39__50_, u5_mult_82_CARRYB_39__51_,
         u5_mult_82_CARRYB_40__0_, u5_mult_82_CARRYB_40__1_,
         u5_mult_82_CARRYB_40__2_, u5_mult_82_CARRYB_40__3_,
         u5_mult_82_CARRYB_40__4_, u5_mult_82_CARRYB_40__5_,
         u5_mult_82_CARRYB_40__6_, u5_mult_82_CARRYB_40__7_,
         u5_mult_82_CARRYB_40__8_, u5_mult_82_CARRYB_40__9_,
         u5_mult_82_CARRYB_40__10_, u5_mult_82_CARRYB_40__11_,
         u5_mult_82_CARRYB_40__12_, u5_mult_82_CARRYB_40__13_,
         u5_mult_82_CARRYB_40__14_, u5_mult_82_CARRYB_40__15_,
         u5_mult_82_CARRYB_40__16_, u5_mult_82_CARRYB_40__17_,
         u5_mult_82_CARRYB_40__18_, u5_mult_82_CARRYB_40__19_,
         u5_mult_82_CARRYB_40__20_, u5_mult_82_CARRYB_40__21_,
         u5_mult_82_CARRYB_40__22_, u5_mult_82_CARRYB_40__23_,
         u5_mult_82_CARRYB_40__24_, u5_mult_82_CARRYB_40__25_,
         u5_mult_82_CARRYB_40__26_, u5_mult_82_CARRYB_40__27_,
         u5_mult_82_CARRYB_40__28_, u5_mult_82_CARRYB_40__29_,
         u5_mult_82_CARRYB_40__30_, u5_mult_82_CARRYB_40__31_,
         u5_mult_82_CARRYB_40__32_, u5_mult_82_CARRYB_40__33_,
         u5_mult_82_CARRYB_40__34_, u5_mult_82_CARRYB_40__35_,
         u5_mult_82_CARRYB_40__36_, u5_mult_82_CARRYB_40__37_,
         u5_mult_82_CARRYB_40__38_, u5_mult_82_CARRYB_40__39_,
         u5_mult_82_CARRYB_40__40_, u5_mult_82_CARRYB_40__41_,
         u5_mult_82_CARRYB_40__42_, u5_mult_82_CARRYB_40__43_,
         u5_mult_82_CARRYB_40__44_, u5_mult_82_CARRYB_40__45_,
         u5_mult_82_CARRYB_40__46_, u5_mult_82_CARRYB_40__47_,
         u5_mult_82_CARRYB_40__48_, u5_mult_82_CARRYB_40__49_,
         u5_mult_82_CARRYB_40__50_, u5_mult_82_CARRYB_40__51_,
         u5_mult_82_CARRYB_41__0_, u5_mult_82_CARRYB_41__1_,
         u5_mult_82_CARRYB_41__2_, u5_mult_82_CARRYB_41__3_,
         u5_mult_82_CARRYB_41__4_, u5_mult_82_CARRYB_41__5_,
         u5_mult_82_CARRYB_41__6_, u5_mult_82_CARRYB_41__7_,
         u5_mult_82_CARRYB_41__8_, u5_mult_82_CARRYB_41__9_,
         u5_mult_82_CARRYB_41__10_, u5_mult_82_CARRYB_41__11_,
         u5_mult_82_CARRYB_41__12_, u5_mult_82_CARRYB_41__13_,
         u5_mult_82_CARRYB_41__14_, u5_mult_82_CARRYB_41__15_,
         u5_mult_82_CARRYB_41__16_, u5_mult_82_CARRYB_41__17_,
         u5_mult_82_CARRYB_41__18_, u5_mult_82_CARRYB_41__19_,
         u5_mult_82_CARRYB_41__20_, u5_mult_82_CARRYB_41__21_,
         u5_mult_82_CARRYB_41__22_, u5_mult_82_CARRYB_41__23_,
         u5_mult_82_CARRYB_41__24_, u5_mult_82_CARRYB_41__25_,
         u5_mult_82_CARRYB_41__26_, u5_mult_82_CARRYB_41__27_,
         u5_mult_82_CARRYB_41__28_, u5_mult_82_CARRYB_41__29_,
         u5_mult_82_CARRYB_41__30_, u5_mult_82_CARRYB_41__31_,
         u5_mult_82_CARRYB_41__32_, u5_mult_82_CARRYB_41__33_,
         u5_mult_82_CARRYB_41__34_, u5_mult_82_CARRYB_41__35_,
         u5_mult_82_CARRYB_41__36_, u5_mult_82_CARRYB_41__37_,
         u5_mult_82_CARRYB_41__38_, u5_mult_82_CARRYB_41__39_,
         u5_mult_82_CARRYB_41__40_, u5_mult_82_CARRYB_41__41_,
         u5_mult_82_CARRYB_41__42_, u5_mult_82_CARRYB_41__43_,
         u5_mult_82_CARRYB_41__44_, u5_mult_82_CARRYB_41__45_,
         u5_mult_82_CARRYB_41__46_, u5_mult_82_CARRYB_41__47_,
         u5_mult_82_CARRYB_41__48_, u5_mult_82_CARRYB_41__49_,
         u5_mult_82_CARRYB_41__50_, u5_mult_82_CARRYB_41__51_,
         u5_mult_82_CARRYB_42__0_, u5_mult_82_CARRYB_42__1_,
         u5_mult_82_CARRYB_42__2_, u5_mult_82_CARRYB_42__3_,
         u5_mult_82_CARRYB_42__4_, u5_mult_82_CARRYB_42__5_,
         u5_mult_82_CARRYB_42__6_, u5_mult_82_CARRYB_42__7_,
         u5_mult_82_CARRYB_42__8_, u5_mult_82_CARRYB_42__9_,
         u5_mult_82_CARRYB_42__10_, u5_mult_82_CARRYB_42__11_,
         u5_mult_82_CARRYB_42__12_, u5_mult_82_CARRYB_42__13_,
         u5_mult_82_CARRYB_42__14_, u5_mult_82_CARRYB_42__15_,
         u5_mult_82_CARRYB_42__16_, u5_mult_82_CARRYB_42__17_,
         u5_mult_82_CARRYB_42__18_, u5_mult_82_CARRYB_42__19_,
         u5_mult_82_CARRYB_42__20_, u5_mult_82_CARRYB_42__21_,
         u5_mult_82_CARRYB_42__22_, u5_mult_82_CARRYB_42__23_,
         u5_mult_82_CARRYB_42__24_, u5_mult_82_CARRYB_42__25_,
         u5_mult_82_CARRYB_42__26_, u5_mult_82_CARRYB_42__27_,
         u5_mult_82_CARRYB_42__28_, u5_mult_82_CARRYB_42__29_,
         u5_mult_82_CARRYB_42__30_, u5_mult_82_CARRYB_42__31_,
         u5_mult_82_CARRYB_42__32_, u5_mult_82_CARRYB_42__33_,
         u5_mult_82_CARRYB_42__34_, u5_mult_82_CARRYB_42__35_,
         u5_mult_82_CARRYB_42__36_, u5_mult_82_CARRYB_42__37_,
         u5_mult_82_CARRYB_42__38_, u5_mult_82_CARRYB_42__39_,
         u5_mult_82_CARRYB_42__40_, u5_mult_82_CARRYB_42__41_,
         u5_mult_82_CARRYB_42__42_, u5_mult_82_CARRYB_42__43_,
         u5_mult_82_CARRYB_42__44_, u5_mult_82_CARRYB_42__45_,
         u5_mult_82_CARRYB_42__46_, u5_mult_82_CARRYB_42__47_,
         u5_mult_82_CARRYB_42__48_, u5_mult_82_CARRYB_42__49_,
         u5_mult_82_CARRYB_42__50_, u5_mult_82_CARRYB_42__51_,
         u5_mult_82_CARRYB_43__0_, u5_mult_82_CARRYB_43__1_,
         u5_mult_82_CARRYB_43__2_, u5_mult_82_CARRYB_43__3_,
         u5_mult_82_CARRYB_43__4_, u5_mult_82_CARRYB_43__5_,
         u5_mult_82_CARRYB_43__6_, u5_mult_82_CARRYB_43__7_,
         u5_mult_82_CARRYB_43__8_, u5_mult_82_CARRYB_43__9_,
         u5_mult_82_CARRYB_43__10_, u5_mult_82_CARRYB_43__11_,
         u5_mult_82_CARRYB_43__12_, u5_mult_82_CARRYB_43__13_,
         u5_mult_82_CARRYB_43__14_, u5_mult_82_CARRYB_43__15_,
         u5_mult_82_CARRYB_43__16_, u5_mult_82_CARRYB_43__17_,
         u5_mult_82_SUMB_24__1_, u5_mult_82_SUMB_24__2_,
         u5_mult_82_SUMB_24__3_, u5_mult_82_SUMB_24__4_,
         u5_mult_82_SUMB_24__5_, u5_mult_82_SUMB_24__6_,
         u5_mult_82_SUMB_24__7_, u5_mult_82_SUMB_24__8_,
         u5_mult_82_SUMB_24__9_, u5_mult_82_SUMB_24__10_,
         u5_mult_82_SUMB_24__11_, u5_mult_82_SUMB_24__12_,
         u5_mult_82_SUMB_24__13_, u5_mult_82_SUMB_24__14_,
         u5_mult_82_SUMB_24__15_, u5_mult_82_SUMB_24__16_,
         u5_mult_82_SUMB_24__17_, u5_mult_82_SUMB_24__18_,
         u5_mult_82_SUMB_24__19_, u5_mult_82_SUMB_24__20_,
         u5_mult_82_SUMB_24__21_, u5_mult_82_SUMB_24__22_,
         u5_mult_82_SUMB_24__23_, u5_mult_82_SUMB_24__24_,
         u5_mult_82_SUMB_24__25_, u5_mult_82_SUMB_24__26_,
         u5_mult_82_SUMB_24__27_, u5_mult_82_SUMB_24__28_,
         u5_mult_82_SUMB_24__29_, u5_mult_82_SUMB_24__30_,
         u5_mult_82_SUMB_24__31_, u5_mult_82_SUMB_24__32_,
         u5_mult_82_SUMB_24__33_, u5_mult_82_SUMB_24__34_,
         u5_mult_82_SUMB_24__35_, u5_mult_82_SUMB_24__36_,
         u5_mult_82_SUMB_24__37_, u5_mult_82_SUMB_24__38_,
         u5_mult_82_SUMB_24__39_, u5_mult_82_SUMB_24__40_,
         u5_mult_82_SUMB_24__41_, u5_mult_82_SUMB_24__42_,
         u5_mult_82_SUMB_24__43_, u5_mult_82_SUMB_24__44_,
         u5_mult_82_SUMB_24__45_, u5_mult_82_SUMB_24__46_,
         u5_mult_82_SUMB_24__47_, u5_mult_82_SUMB_24__48_,
         u5_mult_82_SUMB_24__49_, u5_mult_82_SUMB_24__50_,
         u5_mult_82_SUMB_24__51_, u5_mult_82_SUMB_25__1_,
         u5_mult_82_SUMB_25__2_, u5_mult_82_SUMB_25__3_,
         u5_mult_82_SUMB_25__4_, u5_mult_82_SUMB_25__5_,
         u5_mult_82_SUMB_25__6_, u5_mult_82_SUMB_25__7_,
         u5_mult_82_SUMB_25__8_, u5_mult_82_SUMB_25__9_,
         u5_mult_82_SUMB_25__10_, u5_mult_82_SUMB_25__11_,
         u5_mult_82_SUMB_25__12_, u5_mult_82_SUMB_25__13_,
         u5_mult_82_SUMB_25__14_, u5_mult_82_SUMB_25__15_,
         u5_mult_82_SUMB_25__16_, u5_mult_82_SUMB_25__17_,
         u5_mult_82_SUMB_25__18_, u5_mult_82_SUMB_25__19_,
         u5_mult_82_SUMB_25__20_, u5_mult_82_SUMB_25__21_,
         u5_mult_82_SUMB_25__22_, u5_mult_82_SUMB_25__23_,
         u5_mult_82_SUMB_25__24_, u5_mult_82_SUMB_25__25_,
         u5_mult_82_SUMB_25__26_, u5_mult_82_SUMB_25__27_,
         u5_mult_82_SUMB_25__28_, u5_mult_82_SUMB_25__29_,
         u5_mult_82_SUMB_25__30_, u5_mult_82_SUMB_25__31_,
         u5_mult_82_SUMB_25__32_, u5_mult_82_SUMB_25__33_,
         u5_mult_82_SUMB_25__34_, u5_mult_82_SUMB_25__35_,
         u5_mult_82_SUMB_25__36_, u5_mult_82_SUMB_25__37_,
         u5_mult_82_SUMB_25__38_, u5_mult_82_SUMB_25__39_,
         u5_mult_82_SUMB_25__40_, u5_mult_82_SUMB_25__41_,
         u5_mult_82_SUMB_25__42_, u5_mult_82_SUMB_25__43_,
         u5_mult_82_SUMB_25__44_, u5_mult_82_SUMB_25__45_,
         u5_mult_82_SUMB_25__46_, u5_mult_82_SUMB_25__47_,
         u5_mult_82_SUMB_25__48_, u5_mult_82_SUMB_25__49_,
         u5_mult_82_SUMB_25__50_, u5_mult_82_SUMB_25__51_,
         u5_mult_82_SUMB_26__1_, u5_mult_82_SUMB_26__2_,
         u5_mult_82_SUMB_26__3_, u5_mult_82_SUMB_26__4_,
         u5_mult_82_SUMB_26__5_, u5_mult_82_SUMB_26__6_,
         u5_mult_82_SUMB_26__7_, u5_mult_82_SUMB_26__8_,
         u5_mult_82_SUMB_26__9_, u5_mult_82_SUMB_26__10_,
         u5_mult_82_SUMB_26__11_, u5_mult_82_SUMB_26__12_,
         u5_mult_82_SUMB_26__13_, u5_mult_82_SUMB_26__14_,
         u5_mult_82_SUMB_26__15_, u5_mult_82_SUMB_26__16_,
         u5_mult_82_SUMB_26__17_, u5_mult_82_SUMB_26__18_,
         u5_mult_82_SUMB_26__19_, u5_mult_82_SUMB_26__20_,
         u5_mult_82_SUMB_26__21_, u5_mult_82_SUMB_26__22_,
         u5_mult_82_SUMB_26__23_, u5_mult_82_SUMB_26__24_,
         u5_mult_82_SUMB_26__25_, u5_mult_82_SUMB_26__26_,
         u5_mult_82_SUMB_26__27_, u5_mult_82_SUMB_26__28_,
         u5_mult_82_SUMB_26__29_, u5_mult_82_SUMB_26__30_,
         u5_mult_82_SUMB_26__31_, u5_mult_82_SUMB_26__32_,
         u5_mult_82_SUMB_26__33_, u5_mult_82_SUMB_26__34_,
         u5_mult_82_SUMB_26__35_, u5_mult_82_SUMB_26__36_,
         u5_mult_82_SUMB_26__37_, u5_mult_82_SUMB_26__38_,
         u5_mult_82_SUMB_26__39_, u5_mult_82_SUMB_26__40_,
         u5_mult_82_SUMB_26__41_, u5_mult_82_SUMB_26__42_,
         u5_mult_82_SUMB_26__43_, u5_mult_82_SUMB_26__44_,
         u5_mult_82_SUMB_26__45_, u5_mult_82_SUMB_26__46_,
         u5_mult_82_SUMB_26__47_, u5_mult_82_SUMB_26__48_,
         u5_mult_82_SUMB_26__49_, u5_mult_82_SUMB_26__50_,
         u5_mult_82_SUMB_26__51_, u5_mult_82_SUMB_27__1_,
         u5_mult_82_SUMB_27__2_, u5_mult_82_SUMB_27__3_,
         u5_mult_82_SUMB_27__4_, u5_mult_82_SUMB_27__5_,
         u5_mult_82_SUMB_27__6_, u5_mult_82_SUMB_27__7_,
         u5_mult_82_SUMB_27__8_, u5_mult_82_SUMB_27__9_,
         u5_mult_82_SUMB_27__10_, u5_mult_82_SUMB_27__11_,
         u5_mult_82_SUMB_27__12_, u5_mult_82_SUMB_27__13_,
         u5_mult_82_SUMB_27__14_, u5_mult_82_SUMB_27__15_,
         u5_mult_82_SUMB_27__16_, u5_mult_82_SUMB_27__17_,
         u5_mult_82_SUMB_27__18_, u5_mult_82_SUMB_27__19_,
         u5_mult_82_SUMB_27__20_, u5_mult_82_SUMB_27__21_,
         u5_mult_82_SUMB_27__22_, u5_mult_82_SUMB_27__23_,
         u5_mult_82_SUMB_27__24_, u5_mult_82_SUMB_27__25_,
         u5_mult_82_SUMB_27__26_, u5_mult_82_SUMB_27__27_,
         u5_mult_82_SUMB_27__28_, u5_mult_82_SUMB_27__29_,
         u5_mult_82_SUMB_27__30_, u5_mult_82_SUMB_27__31_,
         u5_mult_82_SUMB_27__32_, u5_mult_82_SUMB_27__33_,
         u5_mult_82_SUMB_27__34_, u5_mult_82_SUMB_27__35_,
         u5_mult_82_SUMB_27__36_, u5_mult_82_SUMB_27__37_,
         u5_mult_82_SUMB_27__38_, u5_mult_82_SUMB_27__39_,
         u5_mult_82_SUMB_27__40_, u5_mult_82_SUMB_27__41_,
         u5_mult_82_SUMB_27__42_, u5_mult_82_SUMB_27__43_,
         u5_mult_82_SUMB_27__44_, u5_mult_82_SUMB_27__45_,
         u5_mult_82_SUMB_27__46_, u5_mult_82_SUMB_27__47_,
         u5_mult_82_SUMB_27__48_, u5_mult_82_SUMB_27__49_,
         u5_mult_82_SUMB_27__50_, u5_mult_82_SUMB_27__51_,
         u5_mult_82_SUMB_28__1_, u5_mult_82_SUMB_28__2_,
         u5_mult_82_SUMB_28__3_, u5_mult_82_SUMB_28__4_,
         u5_mult_82_SUMB_28__5_, u5_mult_82_SUMB_28__6_,
         u5_mult_82_SUMB_28__7_, u5_mult_82_SUMB_28__8_,
         u5_mult_82_SUMB_28__9_, u5_mult_82_SUMB_28__10_,
         u5_mult_82_SUMB_28__11_, u5_mult_82_SUMB_28__12_,
         u5_mult_82_SUMB_28__13_, u5_mult_82_SUMB_28__14_,
         u5_mult_82_SUMB_28__15_, u5_mult_82_SUMB_28__16_,
         u5_mult_82_SUMB_28__17_, u5_mult_82_SUMB_28__18_,
         u5_mult_82_SUMB_28__19_, u5_mult_82_SUMB_28__20_,
         u5_mult_82_SUMB_28__21_, u5_mult_82_SUMB_28__22_,
         u5_mult_82_SUMB_28__23_, u5_mult_82_SUMB_28__24_,
         u5_mult_82_SUMB_28__25_, u5_mult_82_SUMB_28__26_,
         u5_mult_82_SUMB_28__27_, u5_mult_82_SUMB_28__28_,
         u5_mult_82_SUMB_28__29_, u5_mult_82_SUMB_28__30_,
         u5_mult_82_SUMB_28__31_, u5_mult_82_SUMB_28__32_,
         u5_mult_82_SUMB_28__33_, u5_mult_82_SUMB_28__34_,
         u5_mult_82_SUMB_28__35_, u5_mult_82_SUMB_28__36_,
         u5_mult_82_SUMB_28__37_, u5_mult_82_SUMB_28__38_,
         u5_mult_82_SUMB_28__39_, u5_mult_82_SUMB_28__40_,
         u5_mult_82_SUMB_28__41_, u5_mult_82_SUMB_28__42_,
         u5_mult_82_SUMB_28__43_, u5_mult_82_SUMB_28__44_,
         u5_mult_82_SUMB_28__45_, u5_mult_82_SUMB_28__46_,
         u5_mult_82_SUMB_28__47_, u5_mult_82_SUMB_28__48_,
         u5_mult_82_SUMB_28__49_, u5_mult_82_SUMB_28__50_,
         u5_mult_82_SUMB_28__51_, u5_mult_82_SUMB_29__1_,
         u5_mult_82_SUMB_29__2_, u5_mult_82_SUMB_29__3_,
         u5_mult_82_SUMB_29__4_, u5_mult_82_SUMB_29__5_,
         u5_mult_82_SUMB_29__6_, u5_mult_82_SUMB_29__7_,
         u5_mult_82_SUMB_29__8_, u5_mult_82_SUMB_29__9_,
         u5_mult_82_SUMB_29__10_, u5_mult_82_SUMB_29__11_,
         u5_mult_82_SUMB_29__12_, u5_mult_82_SUMB_29__13_,
         u5_mult_82_SUMB_29__14_, u5_mult_82_SUMB_29__15_,
         u5_mult_82_SUMB_29__16_, u5_mult_82_SUMB_29__17_,
         u5_mult_82_SUMB_29__18_, u5_mult_82_SUMB_29__19_,
         u5_mult_82_SUMB_29__20_, u5_mult_82_SUMB_29__21_,
         u5_mult_82_SUMB_29__22_, u5_mult_82_SUMB_29__23_,
         u5_mult_82_SUMB_29__24_, u5_mult_82_SUMB_29__25_,
         u5_mult_82_SUMB_29__26_, u5_mult_82_SUMB_29__27_,
         u5_mult_82_SUMB_29__28_, u5_mult_82_SUMB_29__29_,
         u5_mult_82_SUMB_29__30_, u5_mult_82_SUMB_29__31_,
         u5_mult_82_SUMB_29__32_, u5_mult_82_SUMB_29__33_,
         u5_mult_82_SUMB_29__34_, u5_mult_82_SUMB_29__35_,
         u5_mult_82_SUMB_29__36_, u5_mult_82_SUMB_29__37_,
         u5_mult_82_SUMB_29__38_, u5_mult_82_SUMB_29__39_,
         u5_mult_82_SUMB_29__40_, u5_mult_82_SUMB_29__41_,
         u5_mult_82_SUMB_29__42_, u5_mult_82_SUMB_29__43_,
         u5_mult_82_SUMB_29__44_, u5_mult_82_SUMB_29__45_,
         u5_mult_82_SUMB_29__46_, u5_mult_82_SUMB_29__47_,
         u5_mult_82_SUMB_29__48_, u5_mult_82_SUMB_29__49_,
         u5_mult_82_SUMB_29__50_, u5_mult_82_SUMB_29__51_,
         u5_mult_82_SUMB_30__1_, u5_mult_82_SUMB_30__2_,
         u5_mult_82_SUMB_30__3_, u5_mult_82_SUMB_30__4_,
         u5_mult_82_SUMB_30__5_, u5_mult_82_SUMB_30__6_,
         u5_mult_82_SUMB_30__7_, u5_mult_82_SUMB_30__8_,
         u5_mult_82_SUMB_30__9_, u5_mult_82_SUMB_30__10_,
         u5_mult_82_SUMB_30__11_, u5_mult_82_SUMB_30__12_,
         u5_mult_82_SUMB_30__13_, u5_mult_82_SUMB_30__14_,
         u5_mult_82_SUMB_30__15_, u5_mult_82_SUMB_30__16_,
         u5_mult_82_SUMB_30__17_, u5_mult_82_SUMB_30__18_,
         u5_mult_82_SUMB_30__19_, u5_mult_82_SUMB_30__20_,
         u5_mult_82_SUMB_30__21_, u5_mult_82_SUMB_30__22_,
         u5_mult_82_SUMB_30__23_, u5_mult_82_SUMB_30__24_,
         u5_mult_82_SUMB_30__25_, u5_mult_82_SUMB_30__26_,
         u5_mult_82_SUMB_30__27_, u5_mult_82_SUMB_30__28_,
         u5_mult_82_SUMB_30__29_, u5_mult_82_SUMB_30__30_,
         u5_mult_82_SUMB_30__31_, u5_mult_82_SUMB_30__32_,
         u5_mult_82_SUMB_30__33_, u5_mult_82_SUMB_30__34_,
         u5_mult_82_SUMB_30__35_, u5_mult_82_SUMB_30__36_,
         u5_mult_82_SUMB_30__37_, u5_mult_82_SUMB_30__38_,
         u5_mult_82_SUMB_30__39_, u5_mult_82_SUMB_30__40_,
         u5_mult_82_SUMB_30__41_, u5_mult_82_SUMB_30__42_,
         u5_mult_82_SUMB_30__43_, u5_mult_82_SUMB_30__44_,
         u5_mult_82_SUMB_30__45_, u5_mult_82_SUMB_30__46_,
         u5_mult_82_SUMB_30__47_, u5_mult_82_SUMB_30__48_,
         u5_mult_82_SUMB_30__49_, u5_mult_82_SUMB_30__50_,
         u5_mult_82_SUMB_30__51_, u5_mult_82_SUMB_31__1_,
         u5_mult_82_SUMB_31__2_, u5_mult_82_SUMB_31__3_,
         u5_mult_82_SUMB_31__4_, u5_mult_82_SUMB_31__5_,
         u5_mult_82_SUMB_31__6_, u5_mult_82_SUMB_31__7_,
         u5_mult_82_SUMB_31__8_, u5_mult_82_SUMB_31__9_,
         u5_mult_82_SUMB_31__10_, u5_mult_82_SUMB_31__11_,
         u5_mult_82_SUMB_31__12_, u5_mult_82_SUMB_31__13_,
         u5_mult_82_SUMB_31__14_, u5_mult_82_SUMB_31__15_,
         u5_mult_82_SUMB_31__16_, u5_mult_82_SUMB_31__17_,
         u5_mult_82_SUMB_31__18_, u5_mult_82_SUMB_31__19_,
         u5_mult_82_SUMB_31__20_, u5_mult_82_SUMB_31__21_,
         u5_mult_82_SUMB_31__22_, u5_mult_82_SUMB_31__23_,
         u5_mult_82_SUMB_31__24_, u5_mult_82_SUMB_31__25_,
         u5_mult_82_SUMB_31__26_, u5_mult_82_SUMB_31__27_,
         u5_mult_82_SUMB_31__28_, u5_mult_82_SUMB_31__29_,
         u5_mult_82_SUMB_31__30_, u5_mult_82_SUMB_31__31_,
         u5_mult_82_SUMB_31__32_, u5_mult_82_SUMB_31__33_,
         u5_mult_82_SUMB_31__34_, u5_mult_82_SUMB_31__35_,
         u5_mult_82_SUMB_31__36_, u5_mult_82_SUMB_31__37_,
         u5_mult_82_SUMB_31__38_, u5_mult_82_SUMB_31__39_,
         u5_mult_82_SUMB_31__40_, u5_mult_82_SUMB_31__41_,
         u5_mult_82_SUMB_31__42_, u5_mult_82_SUMB_31__43_,
         u5_mult_82_SUMB_31__44_, u5_mult_82_SUMB_31__45_,
         u5_mult_82_SUMB_31__46_, u5_mult_82_SUMB_31__47_,
         u5_mult_82_SUMB_31__48_, u5_mult_82_SUMB_31__49_,
         u5_mult_82_SUMB_31__50_, u5_mult_82_SUMB_31__51_,
         u5_mult_82_SUMB_32__1_, u5_mult_82_SUMB_32__2_,
         u5_mult_82_SUMB_32__3_, u5_mult_82_SUMB_32__4_,
         u5_mult_82_SUMB_32__5_, u5_mult_82_SUMB_32__6_,
         u5_mult_82_SUMB_32__7_, u5_mult_82_SUMB_32__8_,
         u5_mult_82_SUMB_32__9_, u5_mult_82_SUMB_32__10_,
         u5_mult_82_SUMB_32__11_, u5_mult_82_SUMB_32__12_,
         u5_mult_82_SUMB_32__13_, u5_mult_82_SUMB_32__14_,
         u5_mult_82_SUMB_32__15_, u5_mult_82_SUMB_32__16_,
         u5_mult_82_SUMB_32__17_, u5_mult_82_SUMB_32__18_,
         u5_mult_82_SUMB_32__19_, u5_mult_82_SUMB_32__20_,
         u5_mult_82_SUMB_32__21_, u5_mult_82_SUMB_32__22_,
         u5_mult_82_SUMB_32__23_, u5_mult_82_SUMB_32__24_,
         u5_mult_82_SUMB_32__25_, u5_mult_82_SUMB_32__26_,
         u5_mult_82_SUMB_32__27_, u5_mult_82_SUMB_32__28_,
         u5_mult_82_SUMB_32__29_, u5_mult_82_SUMB_32__30_,
         u5_mult_82_SUMB_32__31_, u5_mult_82_SUMB_32__32_,
         u5_mult_82_SUMB_32__33_, u5_mult_82_SUMB_32__34_,
         u5_mult_82_SUMB_32__35_, u5_mult_82_SUMB_32__36_,
         u5_mult_82_SUMB_32__37_, u5_mult_82_SUMB_32__38_,
         u5_mult_82_SUMB_32__39_, u5_mult_82_SUMB_32__40_,
         u5_mult_82_SUMB_32__41_, u5_mult_82_SUMB_32__42_,
         u5_mult_82_SUMB_32__43_, u5_mult_82_SUMB_32__44_,
         u5_mult_82_SUMB_32__45_, u5_mult_82_SUMB_32__46_,
         u5_mult_82_SUMB_32__47_, u5_mult_82_SUMB_32__48_,
         u5_mult_82_SUMB_32__49_, u5_mult_82_SUMB_32__50_,
         u5_mult_82_SUMB_32__51_, u5_mult_82_SUMB_33__1_,
         u5_mult_82_SUMB_33__2_, u5_mult_82_SUMB_33__3_,
         u5_mult_82_SUMB_33__4_, u5_mult_82_SUMB_33__5_,
         u5_mult_82_SUMB_33__6_, u5_mult_82_SUMB_33__7_,
         u5_mult_82_SUMB_33__8_, u5_mult_82_SUMB_33__9_,
         u5_mult_82_SUMB_33__10_, u5_mult_82_SUMB_33__11_,
         u5_mult_82_SUMB_33__12_, u5_mult_82_SUMB_33__13_,
         u5_mult_82_SUMB_33__14_, u5_mult_82_SUMB_33__15_,
         u5_mult_82_SUMB_33__16_, u5_mult_82_SUMB_33__17_,
         u5_mult_82_SUMB_33__18_, u5_mult_82_SUMB_33__19_,
         u5_mult_82_SUMB_33__20_, u5_mult_82_SUMB_33__21_,
         u5_mult_82_SUMB_33__22_, u5_mult_82_SUMB_33__23_,
         u5_mult_82_SUMB_33__24_, u5_mult_82_SUMB_33__25_,
         u5_mult_82_SUMB_33__26_, u5_mult_82_SUMB_33__27_,
         u5_mult_82_SUMB_33__28_, u5_mult_82_SUMB_33__29_,
         u5_mult_82_SUMB_33__30_, u5_mult_82_SUMB_33__31_,
         u5_mult_82_SUMB_33__32_, u5_mult_82_SUMB_33__33_,
         u5_mult_82_SUMB_33__34_, u5_mult_82_SUMB_33__35_,
         u5_mult_82_CARRYB_24__1_, u5_mult_82_CARRYB_24__2_,
         u5_mult_82_CARRYB_24__3_, u5_mult_82_CARRYB_24__4_,
         u5_mult_82_CARRYB_24__5_, u5_mult_82_CARRYB_24__6_,
         u5_mult_82_CARRYB_24__7_, u5_mult_82_CARRYB_24__8_,
         u5_mult_82_CARRYB_24__9_, u5_mult_82_CARRYB_24__10_,
         u5_mult_82_CARRYB_24__11_, u5_mult_82_CARRYB_24__12_,
         u5_mult_82_CARRYB_24__13_, u5_mult_82_CARRYB_24__14_,
         u5_mult_82_CARRYB_24__15_, u5_mult_82_CARRYB_24__16_,
         u5_mult_82_CARRYB_24__17_, u5_mult_82_CARRYB_24__18_,
         u5_mult_82_CARRYB_24__19_, u5_mult_82_CARRYB_24__20_,
         u5_mult_82_CARRYB_24__21_, u5_mult_82_CARRYB_24__22_,
         u5_mult_82_CARRYB_24__23_, u5_mult_82_CARRYB_24__24_,
         u5_mult_82_CARRYB_24__25_, u5_mult_82_CARRYB_24__26_,
         u5_mult_82_CARRYB_24__27_, u5_mult_82_CARRYB_24__28_,
         u5_mult_82_CARRYB_24__29_, u5_mult_82_CARRYB_24__30_,
         u5_mult_82_CARRYB_24__31_, u5_mult_82_CARRYB_24__32_,
         u5_mult_82_CARRYB_24__33_, u5_mult_82_CARRYB_24__34_,
         u5_mult_82_CARRYB_24__35_, u5_mult_82_CARRYB_24__36_,
         u5_mult_82_CARRYB_24__37_, u5_mult_82_CARRYB_24__38_,
         u5_mult_82_CARRYB_24__39_, u5_mult_82_CARRYB_24__40_,
         u5_mult_82_CARRYB_24__41_, u5_mult_82_CARRYB_24__42_,
         u5_mult_82_CARRYB_24__43_, u5_mult_82_CARRYB_24__44_,
         u5_mult_82_CARRYB_24__45_, u5_mult_82_CARRYB_24__46_,
         u5_mult_82_CARRYB_24__47_, u5_mult_82_CARRYB_24__48_,
         u5_mult_82_CARRYB_24__49_, u5_mult_82_CARRYB_24__50_,
         u5_mult_82_CARRYB_24__51_, u5_mult_82_CARRYB_25__0_,
         u5_mult_82_CARRYB_25__1_, u5_mult_82_CARRYB_25__2_,
         u5_mult_82_CARRYB_25__3_, u5_mult_82_CARRYB_25__4_,
         u5_mult_82_CARRYB_25__5_, u5_mult_82_CARRYB_25__6_,
         u5_mult_82_CARRYB_25__7_, u5_mult_82_CARRYB_25__8_,
         u5_mult_82_CARRYB_25__9_, u5_mult_82_CARRYB_25__10_,
         u5_mult_82_CARRYB_25__11_, u5_mult_82_CARRYB_25__12_,
         u5_mult_82_CARRYB_25__13_, u5_mult_82_CARRYB_25__14_,
         u5_mult_82_CARRYB_25__15_, u5_mult_82_CARRYB_25__16_,
         u5_mult_82_CARRYB_25__17_, u5_mult_82_CARRYB_25__18_,
         u5_mult_82_CARRYB_25__19_, u5_mult_82_CARRYB_25__20_,
         u5_mult_82_CARRYB_25__21_, u5_mult_82_CARRYB_25__22_,
         u5_mult_82_CARRYB_25__23_, u5_mult_82_CARRYB_25__24_,
         u5_mult_82_CARRYB_25__25_, u5_mult_82_CARRYB_25__26_,
         u5_mult_82_CARRYB_25__27_, u5_mult_82_CARRYB_25__28_,
         u5_mult_82_CARRYB_25__29_, u5_mult_82_CARRYB_25__30_,
         u5_mult_82_CARRYB_25__31_, u5_mult_82_CARRYB_25__32_,
         u5_mult_82_CARRYB_25__33_, u5_mult_82_CARRYB_25__34_,
         u5_mult_82_CARRYB_25__35_, u5_mult_82_CARRYB_25__36_,
         u5_mult_82_CARRYB_25__37_, u5_mult_82_CARRYB_25__38_,
         u5_mult_82_CARRYB_25__39_, u5_mult_82_CARRYB_25__40_,
         u5_mult_82_CARRYB_25__41_, u5_mult_82_CARRYB_25__42_,
         u5_mult_82_CARRYB_25__43_, u5_mult_82_CARRYB_25__44_,
         u5_mult_82_CARRYB_25__45_, u5_mult_82_CARRYB_25__46_,
         u5_mult_82_CARRYB_25__47_, u5_mult_82_CARRYB_25__48_,
         u5_mult_82_CARRYB_25__49_, u5_mult_82_CARRYB_25__50_,
         u5_mult_82_CARRYB_25__51_, u5_mult_82_CARRYB_26__0_,
         u5_mult_82_CARRYB_26__1_, u5_mult_82_CARRYB_26__2_,
         u5_mult_82_CARRYB_26__3_, u5_mult_82_CARRYB_26__4_,
         u5_mult_82_CARRYB_26__5_, u5_mult_82_CARRYB_26__6_,
         u5_mult_82_CARRYB_26__7_, u5_mult_82_CARRYB_26__8_,
         u5_mult_82_CARRYB_26__9_, u5_mult_82_CARRYB_26__10_,
         u5_mult_82_CARRYB_26__11_, u5_mult_82_CARRYB_26__12_,
         u5_mult_82_CARRYB_26__13_, u5_mult_82_CARRYB_26__14_,
         u5_mult_82_CARRYB_26__15_, u5_mult_82_CARRYB_26__16_,
         u5_mult_82_CARRYB_26__17_, u5_mult_82_CARRYB_26__18_,
         u5_mult_82_CARRYB_26__19_, u5_mult_82_CARRYB_26__20_,
         u5_mult_82_CARRYB_26__21_, u5_mult_82_CARRYB_26__22_,
         u5_mult_82_CARRYB_26__23_, u5_mult_82_CARRYB_26__24_,
         u5_mult_82_CARRYB_26__25_, u5_mult_82_CARRYB_26__26_,
         u5_mult_82_CARRYB_26__27_, u5_mult_82_CARRYB_26__28_,
         u5_mult_82_CARRYB_26__29_, u5_mult_82_CARRYB_26__30_,
         u5_mult_82_CARRYB_26__31_, u5_mult_82_CARRYB_26__32_,
         u5_mult_82_CARRYB_26__33_, u5_mult_82_CARRYB_26__34_,
         u5_mult_82_CARRYB_26__35_, u5_mult_82_CARRYB_26__36_,
         u5_mult_82_CARRYB_26__37_, u5_mult_82_CARRYB_26__38_,
         u5_mult_82_CARRYB_26__39_, u5_mult_82_CARRYB_26__40_,
         u5_mult_82_CARRYB_26__41_, u5_mult_82_CARRYB_26__42_,
         u5_mult_82_CARRYB_26__43_, u5_mult_82_CARRYB_26__44_,
         u5_mult_82_CARRYB_26__45_, u5_mult_82_CARRYB_26__46_,
         u5_mult_82_CARRYB_26__47_, u5_mult_82_CARRYB_26__48_,
         u5_mult_82_CARRYB_26__49_, u5_mult_82_CARRYB_26__50_,
         u5_mult_82_CARRYB_26__51_, u5_mult_82_CARRYB_27__0_,
         u5_mult_82_CARRYB_27__1_, u5_mult_82_CARRYB_27__2_,
         u5_mult_82_CARRYB_27__3_, u5_mult_82_CARRYB_27__4_,
         u5_mult_82_CARRYB_27__5_, u5_mult_82_CARRYB_27__6_,
         u5_mult_82_CARRYB_27__7_, u5_mult_82_CARRYB_27__8_,
         u5_mult_82_CARRYB_27__9_, u5_mult_82_CARRYB_27__10_,
         u5_mult_82_CARRYB_27__11_, u5_mult_82_CARRYB_27__12_,
         u5_mult_82_CARRYB_27__13_, u5_mult_82_CARRYB_27__14_,
         u5_mult_82_CARRYB_27__15_, u5_mult_82_CARRYB_27__16_,
         u5_mult_82_CARRYB_27__17_, u5_mult_82_CARRYB_27__18_,
         u5_mult_82_CARRYB_27__19_, u5_mult_82_CARRYB_27__20_,
         u5_mult_82_CARRYB_27__21_, u5_mult_82_CARRYB_27__22_,
         u5_mult_82_CARRYB_27__23_, u5_mult_82_CARRYB_27__24_,
         u5_mult_82_CARRYB_27__25_, u5_mult_82_CARRYB_27__26_,
         u5_mult_82_CARRYB_27__27_, u5_mult_82_CARRYB_27__28_,
         u5_mult_82_CARRYB_27__29_, u5_mult_82_CARRYB_27__30_,
         u5_mult_82_CARRYB_27__31_, u5_mult_82_CARRYB_27__32_,
         u5_mult_82_CARRYB_27__33_, u5_mult_82_CARRYB_27__34_,
         u5_mult_82_CARRYB_27__35_, u5_mult_82_CARRYB_27__36_,
         u5_mult_82_CARRYB_27__37_, u5_mult_82_CARRYB_27__38_,
         u5_mult_82_CARRYB_27__39_, u5_mult_82_CARRYB_27__40_,
         u5_mult_82_CARRYB_27__41_, u5_mult_82_CARRYB_27__42_,
         u5_mult_82_CARRYB_27__43_, u5_mult_82_CARRYB_27__44_,
         u5_mult_82_CARRYB_27__45_, u5_mult_82_CARRYB_27__46_,
         u5_mult_82_CARRYB_27__47_, u5_mult_82_CARRYB_27__48_,
         u5_mult_82_CARRYB_27__49_, u5_mult_82_CARRYB_27__50_,
         u5_mult_82_CARRYB_27__51_, u5_mult_82_CARRYB_28__0_,
         u5_mult_82_CARRYB_28__1_, u5_mult_82_CARRYB_28__2_,
         u5_mult_82_CARRYB_28__3_, u5_mult_82_CARRYB_28__4_,
         u5_mult_82_CARRYB_28__5_, u5_mult_82_CARRYB_28__6_,
         u5_mult_82_CARRYB_28__7_, u5_mult_82_CARRYB_28__8_,
         u5_mult_82_CARRYB_28__9_, u5_mult_82_CARRYB_28__10_,
         u5_mult_82_CARRYB_28__11_, u5_mult_82_CARRYB_28__12_,
         u5_mult_82_CARRYB_28__13_, u5_mult_82_CARRYB_28__14_,
         u5_mult_82_CARRYB_28__15_, u5_mult_82_CARRYB_28__16_,
         u5_mult_82_CARRYB_28__17_, u5_mult_82_CARRYB_28__18_,
         u5_mult_82_CARRYB_28__19_, u5_mult_82_CARRYB_28__20_,
         u5_mult_82_CARRYB_28__21_, u5_mult_82_CARRYB_28__22_,
         u5_mult_82_CARRYB_28__23_, u5_mult_82_CARRYB_28__24_,
         u5_mult_82_CARRYB_28__25_, u5_mult_82_CARRYB_28__26_,
         u5_mult_82_CARRYB_28__27_, u5_mult_82_CARRYB_28__28_,
         u5_mult_82_CARRYB_28__29_, u5_mult_82_CARRYB_28__30_,
         u5_mult_82_CARRYB_28__31_, u5_mult_82_CARRYB_28__32_,
         u5_mult_82_CARRYB_28__33_, u5_mult_82_CARRYB_28__34_,
         u5_mult_82_CARRYB_28__35_, u5_mult_82_CARRYB_28__36_,
         u5_mult_82_CARRYB_28__37_, u5_mult_82_CARRYB_28__38_,
         u5_mult_82_CARRYB_28__39_, u5_mult_82_CARRYB_28__40_,
         u5_mult_82_CARRYB_28__41_, u5_mult_82_CARRYB_28__42_,
         u5_mult_82_CARRYB_28__43_, u5_mult_82_CARRYB_28__44_,
         u5_mult_82_CARRYB_28__45_, u5_mult_82_CARRYB_28__46_,
         u5_mult_82_CARRYB_28__47_, u5_mult_82_CARRYB_28__48_,
         u5_mult_82_CARRYB_28__49_, u5_mult_82_CARRYB_28__50_,
         u5_mult_82_CARRYB_28__51_, u5_mult_82_CARRYB_29__0_,
         u5_mult_82_CARRYB_29__1_, u5_mult_82_CARRYB_29__2_,
         u5_mult_82_CARRYB_29__3_, u5_mult_82_CARRYB_29__4_,
         u5_mult_82_CARRYB_29__5_, u5_mult_82_CARRYB_29__6_,
         u5_mult_82_CARRYB_29__7_, u5_mult_82_CARRYB_29__8_,
         u5_mult_82_CARRYB_29__9_, u5_mult_82_CARRYB_29__10_,
         u5_mult_82_CARRYB_29__11_, u5_mult_82_CARRYB_29__12_,
         u5_mult_82_CARRYB_29__13_, u5_mult_82_CARRYB_29__14_,
         u5_mult_82_CARRYB_29__15_, u5_mult_82_CARRYB_29__16_,
         u5_mult_82_CARRYB_29__17_, u5_mult_82_CARRYB_29__18_,
         u5_mult_82_CARRYB_29__19_, u5_mult_82_CARRYB_29__20_,
         u5_mult_82_CARRYB_29__21_, u5_mult_82_CARRYB_29__22_,
         u5_mult_82_CARRYB_29__23_, u5_mult_82_CARRYB_29__24_,
         u5_mult_82_CARRYB_29__25_, u5_mult_82_CARRYB_29__26_,
         u5_mult_82_CARRYB_29__27_, u5_mult_82_CARRYB_29__28_,
         u5_mult_82_CARRYB_29__29_, u5_mult_82_CARRYB_29__30_,
         u5_mult_82_CARRYB_29__31_, u5_mult_82_CARRYB_29__32_,
         u5_mult_82_CARRYB_29__33_, u5_mult_82_CARRYB_29__34_,
         u5_mult_82_CARRYB_29__35_, u5_mult_82_CARRYB_29__36_,
         u5_mult_82_CARRYB_29__37_, u5_mult_82_CARRYB_29__38_,
         u5_mult_82_CARRYB_29__39_, u5_mult_82_CARRYB_29__40_,
         u5_mult_82_CARRYB_29__41_, u5_mult_82_CARRYB_29__42_,
         u5_mult_82_CARRYB_29__43_, u5_mult_82_CARRYB_29__44_,
         u5_mult_82_CARRYB_29__45_, u5_mult_82_CARRYB_29__46_,
         u5_mult_82_CARRYB_29__47_, u5_mult_82_CARRYB_29__48_,
         u5_mult_82_CARRYB_29__49_, u5_mult_82_CARRYB_29__50_,
         u5_mult_82_CARRYB_29__51_, u5_mult_82_CARRYB_30__0_,
         u5_mult_82_CARRYB_30__1_, u5_mult_82_CARRYB_30__2_,
         u5_mult_82_CARRYB_30__3_, u5_mult_82_CARRYB_30__4_,
         u5_mult_82_CARRYB_30__5_, u5_mult_82_CARRYB_30__6_,
         u5_mult_82_CARRYB_30__7_, u5_mult_82_CARRYB_30__8_,
         u5_mult_82_CARRYB_30__9_, u5_mult_82_CARRYB_30__10_,
         u5_mult_82_CARRYB_30__11_, u5_mult_82_CARRYB_30__12_,
         u5_mult_82_CARRYB_30__13_, u5_mult_82_CARRYB_30__14_,
         u5_mult_82_CARRYB_30__15_, u5_mult_82_CARRYB_30__16_,
         u5_mult_82_CARRYB_30__17_, u5_mult_82_CARRYB_30__18_,
         u5_mult_82_CARRYB_30__19_, u5_mult_82_CARRYB_30__20_,
         u5_mult_82_CARRYB_30__21_, u5_mult_82_CARRYB_30__22_,
         u5_mult_82_CARRYB_30__23_, u5_mult_82_CARRYB_30__24_,
         u5_mult_82_CARRYB_30__25_, u5_mult_82_CARRYB_30__26_,
         u5_mult_82_CARRYB_30__27_, u5_mult_82_CARRYB_30__28_,
         u5_mult_82_CARRYB_30__29_, u5_mult_82_CARRYB_30__30_,
         u5_mult_82_CARRYB_30__31_, u5_mult_82_CARRYB_30__32_,
         u5_mult_82_CARRYB_30__33_, u5_mult_82_CARRYB_30__34_,
         u5_mult_82_CARRYB_30__35_, u5_mult_82_CARRYB_30__36_,
         u5_mult_82_CARRYB_30__37_, u5_mult_82_CARRYB_30__38_,
         u5_mult_82_CARRYB_30__39_, u5_mult_82_CARRYB_30__40_,
         u5_mult_82_CARRYB_30__41_, u5_mult_82_CARRYB_30__42_,
         u5_mult_82_CARRYB_30__43_, u5_mult_82_CARRYB_30__44_,
         u5_mult_82_CARRYB_30__45_, u5_mult_82_CARRYB_30__46_,
         u5_mult_82_CARRYB_30__47_, u5_mult_82_CARRYB_30__48_,
         u5_mult_82_CARRYB_30__49_, u5_mult_82_CARRYB_30__50_,
         u5_mult_82_CARRYB_30__51_, u5_mult_82_CARRYB_31__0_,
         u5_mult_82_CARRYB_31__1_, u5_mult_82_CARRYB_31__2_,
         u5_mult_82_CARRYB_31__3_, u5_mult_82_CARRYB_31__4_,
         u5_mult_82_CARRYB_31__5_, u5_mult_82_CARRYB_31__6_,
         u5_mult_82_CARRYB_31__7_, u5_mult_82_CARRYB_31__8_,
         u5_mult_82_CARRYB_31__9_, u5_mult_82_CARRYB_31__10_,
         u5_mult_82_CARRYB_31__11_, u5_mult_82_CARRYB_31__12_,
         u5_mult_82_CARRYB_31__13_, u5_mult_82_CARRYB_31__14_,
         u5_mult_82_CARRYB_31__15_, u5_mult_82_CARRYB_31__16_,
         u5_mult_82_CARRYB_31__17_, u5_mult_82_CARRYB_31__18_,
         u5_mult_82_CARRYB_31__19_, u5_mult_82_CARRYB_31__20_,
         u5_mult_82_CARRYB_31__21_, u5_mult_82_CARRYB_31__22_,
         u5_mult_82_CARRYB_31__23_, u5_mult_82_CARRYB_31__24_,
         u5_mult_82_CARRYB_31__25_, u5_mult_82_CARRYB_31__26_,
         u5_mult_82_CARRYB_31__27_, u5_mult_82_CARRYB_31__28_,
         u5_mult_82_CARRYB_31__29_, u5_mult_82_CARRYB_31__30_,
         u5_mult_82_CARRYB_31__31_, u5_mult_82_CARRYB_31__32_,
         u5_mult_82_CARRYB_31__33_, u5_mult_82_CARRYB_31__34_,
         u5_mult_82_CARRYB_31__35_, u5_mult_82_CARRYB_31__36_,
         u5_mult_82_CARRYB_31__37_, u5_mult_82_CARRYB_31__38_,
         u5_mult_82_CARRYB_31__39_, u5_mult_82_CARRYB_31__40_,
         u5_mult_82_CARRYB_31__41_, u5_mult_82_CARRYB_31__42_,
         u5_mult_82_CARRYB_31__43_, u5_mult_82_CARRYB_31__44_,
         u5_mult_82_CARRYB_31__45_, u5_mult_82_CARRYB_31__46_,
         u5_mult_82_CARRYB_31__47_, u5_mult_82_CARRYB_31__48_,
         u5_mult_82_CARRYB_31__49_, u5_mult_82_CARRYB_31__50_,
         u5_mult_82_CARRYB_31__51_, u5_mult_82_CARRYB_32__0_,
         u5_mult_82_CARRYB_32__1_, u5_mult_82_CARRYB_32__2_,
         u5_mult_82_CARRYB_32__3_, u5_mult_82_CARRYB_32__4_,
         u5_mult_82_CARRYB_32__5_, u5_mult_82_CARRYB_32__6_,
         u5_mult_82_CARRYB_32__7_, u5_mult_82_CARRYB_32__8_,
         u5_mult_82_CARRYB_32__9_, u5_mult_82_CARRYB_32__10_,
         u5_mult_82_CARRYB_32__11_, u5_mult_82_CARRYB_32__12_,
         u5_mult_82_CARRYB_32__13_, u5_mult_82_CARRYB_32__14_,
         u5_mult_82_CARRYB_32__15_, u5_mult_82_CARRYB_32__16_,
         u5_mult_82_CARRYB_32__17_, u5_mult_82_CARRYB_32__18_,
         u5_mult_82_CARRYB_32__19_, u5_mult_82_CARRYB_32__20_,
         u5_mult_82_CARRYB_32__21_, u5_mult_82_CARRYB_32__22_,
         u5_mult_82_CARRYB_32__23_, u5_mult_82_CARRYB_32__24_,
         u5_mult_82_CARRYB_32__25_, u5_mult_82_CARRYB_32__26_,
         u5_mult_82_CARRYB_32__27_, u5_mult_82_CARRYB_32__28_,
         u5_mult_82_CARRYB_32__29_, u5_mult_82_CARRYB_32__30_,
         u5_mult_82_CARRYB_32__31_, u5_mult_82_CARRYB_32__32_,
         u5_mult_82_CARRYB_32__33_, u5_mult_82_CARRYB_32__34_,
         u5_mult_82_CARRYB_32__35_, u5_mult_82_CARRYB_32__36_,
         u5_mult_82_CARRYB_32__37_, u5_mult_82_CARRYB_32__38_,
         u5_mult_82_CARRYB_32__39_, u5_mult_82_CARRYB_32__40_,
         u5_mult_82_CARRYB_32__41_, u5_mult_82_CARRYB_32__42_,
         u5_mult_82_CARRYB_32__43_, u5_mult_82_CARRYB_32__44_,
         u5_mult_82_CARRYB_32__45_, u5_mult_82_CARRYB_32__46_,
         u5_mult_82_CARRYB_32__47_, u5_mult_82_CARRYB_32__48_,
         u5_mult_82_CARRYB_32__49_, u5_mult_82_CARRYB_32__50_,
         u5_mult_82_CARRYB_32__51_, u5_mult_82_CARRYB_33__0_,
         u5_mult_82_CARRYB_33__1_, u5_mult_82_CARRYB_33__2_,
         u5_mult_82_CARRYB_33__3_, u5_mult_82_CARRYB_33__4_,
         u5_mult_82_CARRYB_33__5_, u5_mult_82_CARRYB_33__6_,
         u5_mult_82_CARRYB_33__7_, u5_mult_82_CARRYB_33__8_,
         u5_mult_82_CARRYB_33__9_, u5_mult_82_CARRYB_33__10_,
         u5_mult_82_CARRYB_33__11_, u5_mult_82_CARRYB_33__12_,
         u5_mult_82_CARRYB_33__13_, u5_mult_82_CARRYB_33__14_,
         u5_mult_82_CARRYB_33__15_, u5_mult_82_CARRYB_33__16_,
         u5_mult_82_CARRYB_33__17_, u5_mult_82_CARRYB_33__18_,
         u5_mult_82_CARRYB_33__19_, u5_mult_82_CARRYB_33__20_,
         u5_mult_82_CARRYB_33__21_, u5_mult_82_CARRYB_33__22_,
         u5_mult_82_CARRYB_33__23_, u5_mult_82_CARRYB_33__24_,
         u5_mult_82_CARRYB_33__25_, u5_mult_82_CARRYB_33__26_,
         u5_mult_82_CARRYB_33__27_, u5_mult_82_CARRYB_33__28_,
         u5_mult_82_CARRYB_33__29_, u5_mult_82_CARRYB_33__30_,
         u5_mult_82_CARRYB_33__31_, u5_mult_82_CARRYB_33__32_,
         u5_mult_82_CARRYB_33__33_, u5_mult_82_CARRYB_33__34_,
         u5_mult_82_CARRYB_33__35_, u5_mult_82_SUMB_14__19_,
         u5_mult_82_SUMB_14__20_, u5_mult_82_SUMB_14__21_,
         u5_mult_82_SUMB_14__22_, u5_mult_82_SUMB_14__23_,
         u5_mult_82_SUMB_14__24_, u5_mult_82_SUMB_14__25_,
         u5_mult_82_SUMB_14__26_, u5_mult_82_SUMB_14__27_,
         u5_mult_82_SUMB_14__28_, u5_mult_82_SUMB_14__29_,
         u5_mult_82_SUMB_14__30_, u5_mult_82_SUMB_14__31_,
         u5_mult_82_SUMB_14__32_, u5_mult_82_SUMB_14__33_,
         u5_mult_82_SUMB_14__34_, u5_mult_82_SUMB_14__35_,
         u5_mult_82_SUMB_14__36_, u5_mult_82_SUMB_14__37_,
         u5_mult_82_SUMB_14__38_, u5_mult_82_SUMB_14__39_,
         u5_mult_82_SUMB_14__40_, u5_mult_82_SUMB_14__41_,
         u5_mult_82_SUMB_14__42_, u5_mult_82_SUMB_14__43_,
         u5_mult_82_SUMB_14__44_, u5_mult_82_SUMB_14__45_,
         u5_mult_82_SUMB_14__46_, u5_mult_82_SUMB_14__47_,
         u5_mult_82_SUMB_14__48_, u5_mult_82_SUMB_14__49_,
         u5_mult_82_SUMB_14__50_, u5_mult_82_SUMB_14__51_,
         u5_mult_82_SUMB_15__1_, u5_mult_82_SUMB_15__2_,
         u5_mult_82_SUMB_15__3_, u5_mult_82_SUMB_15__4_,
         u5_mult_82_SUMB_15__5_, u5_mult_82_SUMB_15__6_,
         u5_mult_82_SUMB_15__7_, u5_mult_82_SUMB_15__8_,
         u5_mult_82_SUMB_15__9_, u5_mult_82_SUMB_15__10_,
         u5_mult_82_SUMB_15__11_, u5_mult_82_SUMB_15__12_,
         u5_mult_82_SUMB_15__13_, u5_mult_82_SUMB_15__14_,
         u5_mult_82_SUMB_15__15_, u5_mult_82_SUMB_15__16_,
         u5_mult_82_SUMB_15__17_, u5_mult_82_SUMB_15__18_,
         u5_mult_82_SUMB_15__19_, u5_mult_82_SUMB_15__20_,
         u5_mult_82_SUMB_15__21_, u5_mult_82_SUMB_15__22_,
         u5_mult_82_SUMB_15__23_, u5_mult_82_SUMB_15__24_,
         u5_mult_82_SUMB_15__25_, u5_mult_82_SUMB_15__26_,
         u5_mult_82_SUMB_15__27_, u5_mult_82_SUMB_15__28_,
         u5_mult_82_SUMB_15__29_, u5_mult_82_SUMB_15__30_,
         u5_mult_82_SUMB_15__31_, u5_mult_82_SUMB_15__32_,
         u5_mult_82_SUMB_15__33_, u5_mult_82_SUMB_15__34_,
         u5_mult_82_SUMB_15__35_, u5_mult_82_SUMB_15__36_,
         u5_mult_82_SUMB_15__37_, u5_mult_82_SUMB_15__38_,
         u5_mult_82_SUMB_15__39_, u5_mult_82_SUMB_15__40_,
         u5_mult_82_SUMB_15__41_, u5_mult_82_SUMB_15__42_,
         u5_mult_82_SUMB_15__43_, u5_mult_82_SUMB_15__44_,
         u5_mult_82_SUMB_15__45_, u5_mult_82_SUMB_15__46_,
         u5_mult_82_SUMB_15__47_, u5_mult_82_SUMB_15__48_,
         u5_mult_82_SUMB_15__49_, u5_mult_82_SUMB_15__50_,
         u5_mult_82_SUMB_15__51_, u5_mult_82_SUMB_16__1_,
         u5_mult_82_SUMB_16__2_, u5_mult_82_SUMB_16__3_,
         u5_mult_82_SUMB_16__4_, u5_mult_82_SUMB_16__5_,
         u5_mult_82_SUMB_16__6_, u5_mult_82_SUMB_16__7_,
         u5_mult_82_SUMB_16__8_, u5_mult_82_SUMB_16__9_,
         u5_mult_82_SUMB_16__10_, u5_mult_82_SUMB_16__11_,
         u5_mult_82_SUMB_16__12_, u5_mult_82_SUMB_16__13_,
         u5_mult_82_SUMB_16__14_, u5_mult_82_SUMB_16__15_,
         u5_mult_82_SUMB_16__16_, u5_mult_82_SUMB_16__17_,
         u5_mult_82_SUMB_16__18_, u5_mult_82_SUMB_16__19_,
         u5_mult_82_SUMB_16__20_, u5_mult_82_SUMB_16__21_,
         u5_mult_82_SUMB_16__22_, u5_mult_82_SUMB_16__23_,
         u5_mult_82_SUMB_16__24_, u5_mult_82_SUMB_16__25_,
         u5_mult_82_SUMB_16__26_, u5_mult_82_SUMB_16__27_,
         u5_mult_82_SUMB_16__28_, u5_mult_82_SUMB_16__29_,
         u5_mult_82_SUMB_16__30_, u5_mult_82_SUMB_16__31_,
         u5_mult_82_SUMB_16__32_, u5_mult_82_SUMB_16__33_,
         u5_mult_82_SUMB_16__34_, u5_mult_82_SUMB_16__35_,
         u5_mult_82_SUMB_16__36_, u5_mult_82_SUMB_16__37_,
         u5_mult_82_SUMB_16__38_, u5_mult_82_SUMB_16__39_,
         u5_mult_82_SUMB_16__40_, u5_mult_82_SUMB_16__41_,
         u5_mult_82_SUMB_16__42_, u5_mult_82_SUMB_16__43_,
         u5_mult_82_SUMB_16__44_, u5_mult_82_SUMB_16__45_,
         u5_mult_82_SUMB_16__46_, u5_mult_82_SUMB_16__47_,
         u5_mult_82_SUMB_16__48_, u5_mult_82_SUMB_16__49_,
         u5_mult_82_SUMB_16__50_, u5_mult_82_SUMB_16__51_,
         u5_mult_82_SUMB_17__1_, u5_mult_82_SUMB_17__2_,
         u5_mult_82_SUMB_17__3_, u5_mult_82_SUMB_17__4_,
         u5_mult_82_SUMB_17__5_, u5_mult_82_SUMB_17__6_,
         u5_mult_82_SUMB_17__7_, u5_mult_82_SUMB_17__8_,
         u5_mult_82_SUMB_17__9_, u5_mult_82_SUMB_17__10_,
         u5_mult_82_SUMB_17__11_, u5_mult_82_SUMB_17__12_,
         u5_mult_82_SUMB_17__13_, u5_mult_82_SUMB_17__14_,
         u5_mult_82_SUMB_17__15_, u5_mult_82_SUMB_17__16_,
         u5_mult_82_SUMB_17__17_, u5_mult_82_SUMB_17__18_,
         u5_mult_82_SUMB_17__19_, u5_mult_82_SUMB_17__20_,
         u5_mult_82_SUMB_17__21_, u5_mult_82_SUMB_17__22_,
         u5_mult_82_SUMB_17__23_, u5_mult_82_SUMB_17__24_,
         u5_mult_82_SUMB_17__25_, u5_mult_82_SUMB_17__26_,
         u5_mult_82_SUMB_17__27_, u5_mult_82_SUMB_17__28_,
         u5_mult_82_SUMB_17__29_, u5_mult_82_SUMB_17__30_,
         u5_mult_82_SUMB_17__31_, u5_mult_82_SUMB_17__32_,
         u5_mult_82_SUMB_17__33_, u5_mult_82_SUMB_17__34_,
         u5_mult_82_SUMB_17__35_, u5_mult_82_SUMB_17__36_,
         u5_mult_82_SUMB_17__37_, u5_mult_82_SUMB_17__38_,
         u5_mult_82_SUMB_17__39_, u5_mult_82_SUMB_17__40_,
         u5_mult_82_SUMB_17__41_, u5_mult_82_SUMB_17__42_,
         u5_mult_82_SUMB_17__43_, u5_mult_82_SUMB_17__44_,
         u5_mult_82_SUMB_17__45_, u5_mult_82_SUMB_17__46_,
         u5_mult_82_SUMB_17__47_, u5_mult_82_SUMB_17__48_,
         u5_mult_82_SUMB_17__49_, u5_mult_82_SUMB_17__50_,
         u5_mult_82_SUMB_17__51_, u5_mult_82_SUMB_18__1_,
         u5_mult_82_SUMB_18__2_, u5_mult_82_SUMB_18__3_,
         u5_mult_82_SUMB_18__4_, u5_mult_82_SUMB_18__5_,
         u5_mult_82_SUMB_18__6_, u5_mult_82_SUMB_18__7_,
         u5_mult_82_SUMB_18__8_, u5_mult_82_SUMB_18__9_,
         u5_mult_82_SUMB_18__10_, u5_mult_82_SUMB_18__11_,
         u5_mult_82_SUMB_18__12_, u5_mult_82_SUMB_18__13_,
         u5_mult_82_SUMB_18__14_, u5_mult_82_SUMB_18__15_,
         u5_mult_82_SUMB_18__16_, u5_mult_82_SUMB_18__17_,
         u5_mult_82_SUMB_18__18_, u5_mult_82_SUMB_18__19_,
         u5_mult_82_SUMB_18__20_, u5_mult_82_SUMB_18__21_,
         u5_mult_82_SUMB_18__22_, u5_mult_82_SUMB_18__23_,
         u5_mult_82_SUMB_18__24_, u5_mult_82_SUMB_18__25_,
         u5_mult_82_SUMB_18__26_, u5_mult_82_SUMB_18__27_,
         u5_mult_82_SUMB_18__28_, u5_mult_82_SUMB_18__29_,
         u5_mult_82_SUMB_18__30_, u5_mult_82_SUMB_18__31_,
         u5_mult_82_SUMB_18__32_, u5_mult_82_SUMB_18__33_,
         u5_mult_82_SUMB_18__34_, u5_mult_82_SUMB_18__35_,
         u5_mult_82_SUMB_18__36_, u5_mult_82_SUMB_18__37_,
         u5_mult_82_SUMB_18__38_, u5_mult_82_SUMB_18__39_,
         u5_mult_82_SUMB_18__40_, u5_mult_82_SUMB_18__41_,
         u5_mult_82_SUMB_18__42_, u5_mult_82_SUMB_18__43_,
         u5_mult_82_SUMB_18__44_, u5_mult_82_SUMB_18__45_,
         u5_mult_82_SUMB_18__46_, u5_mult_82_SUMB_18__47_,
         u5_mult_82_SUMB_18__48_, u5_mult_82_SUMB_18__49_,
         u5_mult_82_SUMB_18__50_, u5_mult_82_SUMB_18__51_,
         u5_mult_82_SUMB_19__1_, u5_mult_82_SUMB_19__2_,
         u5_mult_82_SUMB_19__3_, u5_mult_82_SUMB_19__4_,
         u5_mult_82_SUMB_19__5_, u5_mult_82_SUMB_19__6_,
         u5_mult_82_SUMB_19__7_, u5_mult_82_SUMB_19__8_,
         u5_mult_82_SUMB_19__9_, u5_mult_82_SUMB_19__10_,
         u5_mult_82_SUMB_19__11_, u5_mult_82_SUMB_19__12_,
         u5_mult_82_SUMB_19__13_, u5_mult_82_SUMB_19__14_,
         u5_mult_82_SUMB_19__15_, u5_mult_82_SUMB_19__16_,
         u5_mult_82_SUMB_19__17_, u5_mult_82_SUMB_19__18_,
         u5_mult_82_SUMB_19__19_, u5_mult_82_SUMB_19__20_,
         u5_mult_82_SUMB_19__21_, u5_mult_82_SUMB_19__22_,
         u5_mult_82_SUMB_19__23_, u5_mult_82_SUMB_19__24_,
         u5_mult_82_SUMB_19__25_, u5_mult_82_SUMB_19__26_,
         u5_mult_82_SUMB_19__27_, u5_mult_82_SUMB_19__28_,
         u5_mult_82_SUMB_19__29_, u5_mult_82_SUMB_19__30_,
         u5_mult_82_SUMB_19__31_, u5_mult_82_SUMB_19__32_,
         u5_mult_82_SUMB_19__33_, u5_mult_82_SUMB_19__34_,
         u5_mult_82_SUMB_19__35_, u5_mult_82_SUMB_19__36_,
         u5_mult_82_SUMB_19__37_, u5_mult_82_SUMB_19__38_,
         u5_mult_82_SUMB_19__39_, u5_mult_82_SUMB_19__40_,
         u5_mult_82_SUMB_19__41_, u5_mult_82_SUMB_19__42_,
         u5_mult_82_SUMB_19__43_, u5_mult_82_SUMB_19__44_,
         u5_mult_82_SUMB_19__45_, u5_mult_82_SUMB_19__46_,
         u5_mult_82_SUMB_19__47_, u5_mult_82_SUMB_19__48_,
         u5_mult_82_SUMB_19__49_, u5_mult_82_SUMB_19__50_,
         u5_mult_82_SUMB_19__51_, u5_mult_82_SUMB_20__1_,
         u5_mult_82_SUMB_20__2_, u5_mult_82_SUMB_20__3_,
         u5_mult_82_SUMB_20__4_, u5_mult_82_SUMB_20__5_,
         u5_mult_82_SUMB_20__6_, u5_mult_82_SUMB_20__7_,
         u5_mult_82_SUMB_20__8_, u5_mult_82_SUMB_20__9_,
         u5_mult_82_SUMB_20__10_, u5_mult_82_SUMB_20__11_,
         u5_mult_82_SUMB_20__12_, u5_mult_82_SUMB_20__13_,
         u5_mult_82_SUMB_20__14_, u5_mult_82_SUMB_20__15_,
         u5_mult_82_SUMB_20__16_, u5_mult_82_SUMB_20__17_,
         u5_mult_82_SUMB_20__18_, u5_mult_82_SUMB_20__19_,
         u5_mult_82_SUMB_20__20_, u5_mult_82_SUMB_20__21_,
         u5_mult_82_SUMB_20__22_, u5_mult_82_SUMB_20__23_,
         u5_mult_82_SUMB_20__24_, u5_mult_82_SUMB_20__25_,
         u5_mult_82_SUMB_20__26_, u5_mult_82_SUMB_20__27_,
         u5_mult_82_SUMB_20__28_, u5_mult_82_SUMB_20__29_,
         u5_mult_82_SUMB_20__30_, u5_mult_82_SUMB_20__31_,
         u5_mult_82_SUMB_20__32_, u5_mult_82_SUMB_20__33_,
         u5_mult_82_SUMB_20__34_, u5_mult_82_SUMB_20__35_,
         u5_mult_82_SUMB_20__36_, u5_mult_82_SUMB_20__37_,
         u5_mult_82_SUMB_20__38_, u5_mult_82_SUMB_20__39_,
         u5_mult_82_SUMB_20__40_, u5_mult_82_SUMB_20__41_,
         u5_mult_82_SUMB_20__42_, u5_mult_82_SUMB_20__43_,
         u5_mult_82_SUMB_20__44_, u5_mult_82_SUMB_20__45_,
         u5_mult_82_SUMB_20__46_, u5_mult_82_SUMB_20__47_,
         u5_mult_82_SUMB_20__48_, u5_mult_82_SUMB_20__49_,
         u5_mult_82_SUMB_20__50_, u5_mult_82_SUMB_20__51_,
         u5_mult_82_SUMB_21__1_, u5_mult_82_SUMB_21__2_,
         u5_mult_82_SUMB_21__3_, u5_mult_82_SUMB_21__4_,
         u5_mult_82_SUMB_21__5_, u5_mult_82_SUMB_21__6_,
         u5_mult_82_SUMB_21__7_, u5_mult_82_SUMB_21__8_,
         u5_mult_82_SUMB_21__9_, u5_mult_82_SUMB_21__10_,
         u5_mult_82_SUMB_21__11_, u5_mult_82_SUMB_21__12_,
         u5_mult_82_SUMB_21__13_, u5_mult_82_SUMB_21__14_,
         u5_mult_82_SUMB_21__15_, u5_mult_82_SUMB_21__16_,
         u5_mult_82_SUMB_21__17_, u5_mult_82_SUMB_21__18_,
         u5_mult_82_SUMB_21__19_, u5_mult_82_SUMB_21__20_,
         u5_mult_82_SUMB_21__21_, u5_mult_82_SUMB_21__22_,
         u5_mult_82_SUMB_21__23_, u5_mult_82_SUMB_21__24_,
         u5_mult_82_SUMB_21__25_, u5_mult_82_SUMB_21__26_,
         u5_mult_82_SUMB_21__27_, u5_mult_82_SUMB_21__28_,
         u5_mult_82_SUMB_21__29_, u5_mult_82_SUMB_21__30_,
         u5_mult_82_SUMB_21__31_, u5_mult_82_SUMB_21__32_,
         u5_mult_82_SUMB_21__33_, u5_mult_82_SUMB_21__34_,
         u5_mult_82_SUMB_21__35_, u5_mult_82_SUMB_21__36_,
         u5_mult_82_SUMB_21__37_, u5_mult_82_SUMB_21__38_,
         u5_mult_82_SUMB_21__39_, u5_mult_82_SUMB_21__40_,
         u5_mult_82_SUMB_21__41_, u5_mult_82_SUMB_21__42_,
         u5_mult_82_SUMB_21__43_, u5_mult_82_SUMB_21__44_,
         u5_mult_82_SUMB_21__45_, u5_mult_82_SUMB_21__46_,
         u5_mult_82_SUMB_21__47_, u5_mult_82_SUMB_21__48_,
         u5_mult_82_SUMB_21__49_, u5_mult_82_SUMB_21__50_,
         u5_mult_82_SUMB_21__51_, u5_mult_82_SUMB_22__1_,
         u5_mult_82_SUMB_22__2_, u5_mult_82_SUMB_22__3_,
         u5_mult_82_SUMB_22__4_, u5_mult_82_SUMB_22__5_,
         u5_mult_82_SUMB_22__6_, u5_mult_82_SUMB_22__7_,
         u5_mult_82_SUMB_22__8_, u5_mult_82_SUMB_22__9_,
         u5_mult_82_SUMB_22__10_, u5_mult_82_SUMB_22__11_,
         u5_mult_82_SUMB_22__12_, u5_mult_82_SUMB_22__13_,
         u5_mult_82_SUMB_22__14_, u5_mult_82_SUMB_22__15_,
         u5_mult_82_SUMB_22__16_, u5_mult_82_SUMB_22__17_,
         u5_mult_82_SUMB_22__18_, u5_mult_82_SUMB_22__19_,
         u5_mult_82_SUMB_22__20_, u5_mult_82_SUMB_22__21_,
         u5_mult_82_SUMB_22__22_, u5_mult_82_SUMB_22__23_,
         u5_mult_82_SUMB_22__24_, u5_mult_82_SUMB_22__25_,
         u5_mult_82_SUMB_22__26_, u5_mult_82_SUMB_22__27_,
         u5_mult_82_SUMB_22__28_, u5_mult_82_SUMB_22__29_,
         u5_mult_82_SUMB_22__30_, u5_mult_82_SUMB_22__31_,
         u5_mult_82_SUMB_22__32_, u5_mult_82_SUMB_22__33_,
         u5_mult_82_SUMB_22__34_, u5_mult_82_SUMB_22__35_,
         u5_mult_82_SUMB_22__36_, u5_mult_82_SUMB_22__37_,
         u5_mult_82_SUMB_22__38_, u5_mult_82_SUMB_22__39_,
         u5_mult_82_SUMB_22__40_, u5_mult_82_SUMB_22__41_,
         u5_mult_82_SUMB_22__42_, u5_mult_82_SUMB_22__43_,
         u5_mult_82_SUMB_22__44_, u5_mult_82_SUMB_22__45_,
         u5_mult_82_SUMB_22__46_, u5_mult_82_SUMB_22__47_,
         u5_mult_82_SUMB_22__48_, u5_mult_82_SUMB_22__49_,
         u5_mult_82_SUMB_22__50_, u5_mult_82_SUMB_22__51_,
         u5_mult_82_SUMB_23__1_, u5_mult_82_SUMB_23__2_,
         u5_mult_82_SUMB_23__3_, u5_mult_82_SUMB_23__4_,
         u5_mult_82_SUMB_23__5_, u5_mult_82_SUMB_23__6_,
         u5_mult_82_SUMB_23__7_, u5_mult_82_SUMB_23__8_,
         u5_mult_82_SUMB_23__9_, u5_mult_82_SUMB_23__10_,
         u5_mult_82_SUMB_23__11_, u5_mult_82_SUMB_23__12_,
         u5_mult_82_SUMB_23__13_, u5_mult_82_SUMB_23__14_,
         u5_mult_82_SUMB_23__15_, u5_mult_82_SUMB_23__16_,
         u5_mult_82_SUMB_23__17_, u5_mult_82_SUMB_23__18_,
         u5_mult_82_SUMB_23__19_, u5_mult_82_SUMB_23__20_,
         u5_mult_82_SUMB_23__21_, u5_mult_82_SUMB_23__22_,
         u5_mult_82_SUMB_23__23_, u5_mult_82_SUMB_23__24_,
         u5_mult_82_SUMB_23__25_, u5_mult_82_SUMB_23__26_,
         u5_mult_82_SUMB_23__27_, u5_mult_82_SUMB_23__28_,
         u5_mult_82_SUMB_23__29_, u5_mult_82_SUMB_23__30_,
         u5_mult_82_SUMB_23__31_, u5_mult_82_SUMB_23__32_,
         u5_mult_82_SUMB_23__33_, u5_mult_82_SUMB_23__34_,
         u5_mult_82_SUMB_23__35_, u5_mult_82_SUMB_23__36_,
         u5_mult_82_SUMB_23__37_, u5_mult_82_SUMB_23__38_,
         u5_mult_82_SUMB_23__39_, u5_mult_82_SUMB_23__40_,
         u5_mult_82_SUMB_23__41_, u5_mult_82_SUMB_23__42_,
         u5_mult_82_SUMB_23__43_, u5_mult_82_SUMB_23__44_,
         u5_mult_82_SUMB_23__45_, u5_mult_82_SUMB_23__46_,
         u5_mult_82_SUMB_23__47_, u5_mult_82_SUMB_23__48_,
         u5_mult_82_SUMB_23__49_, u5_mult_82_SUMB_23__50_,
         u5_mult_82_SUMB_23__51_, u5_mult_82_CARRYB_14__19_,
         u5_mult_82_CARRYB_14__20_, u5_mult_82_CARRYB_14__21_,
         u5_mult_82_CARRYB_14__22_, u5_mult_82_CARRYB_14__23_,
         u5_mult_82_CARRYB_14__24_, u5_mult_82_CARRYB_14__25_,
         u5_mult_82_CARRYB_14__26_, u5_mult_82_CARRYB_14__27_,
         u5_mult_82_CARRYB_14__28_, u5_mult_82_CARRYB_14__29_,
         u5_mult_82_CARRYB_14__30_, u5_mult_82_CARRYB_14__31_,
         u5_mult_82_CARRYB_14__32_, u5_mult_82_CARRYB_14__33_,
         u5_mult_82_CARRYB_14__34_, u5_mult_82_CARRYB_14__35_,
         u5_mult_82_CARRYB_14__36_, u5_mult_82_CARRYB_14__37_,
         u5_mult_82_CARRYB_14__38_, u5_mult_82_CARRYB_14__39_,
         u5_mult_82_CARRYB_14__40_, u5_mult_82_CARRYB_14__41_,
         u5_mult_82_CARRYB_14__42_, u5_mult_82_CARRYB_14__43_,
         u5_mult_82_CARRYB_14__44_, u5_mult_82_CARRYB_14__45_,
         u5_mult_82_CARRYB_14__46_, u5_mult_82_CARRYB_14__47_,
         u5_mult_82_CARRYB_14__48_, u5_mult_82_CARRYB_14__49_,
         u5_mult_82_CARRYB_14__50_, u5_mult_82_CARRYB_14__51_,
         u5_mult_82_CARRYB_15__0_, u5_mult_82_CARRYB_15__1_,
         u5_mult_82_CARRYB_15__2_, u5_mult_82_CARRYB_15__3_,
         u5_mult_82_CARRYB_15__4_, u5_mult_82_CARRYB_15__5_,
         u5_mult_82_CARRYB_15__6_, u5_mult_82_CARRYB_15__7_,
         u5_mult_82_CARRYB_15__8_, u5_mult_82_CARRYB_15__9_,
         u5_mult_82_CARRYB_15__10_, u5_mult_82_CARRYB_15__11_,
         u5_mult_82_CARRYB_15__12_, u5_mult_82_CARRYB_15__13_,
         u5_mult_82_CARRYB_15__14_, u5_mult_82_CARRYB_15__15_,
         u5_mult_82_CARRYB_15__16_, u5_mult_82_CARRYB_15__17_,
         u5_mult_82_CARRYB_15__18_, u5_mult_82_CARRYB_15__19_,
         u5_mult_82_CARRYB_15__20_, u5_mult_82_CARRYB_15__21_,
         u5_mult_82_CARRYB_15__22_, u5_mult_82_CARRYB_15__23_,
         u5_mult_82_CARRYB_15__24_, u5_mult_82_CARRYB_15__25_,
         u5_mult_82_CARRYB_15__26_, u5_mult_82_CARRYB_15__27_,
         u5_mult_82_CARRYB_15__28_, u5_mult_82_CARRYB_15__29_,
         u5_mult_82_CARRYB_15__30_, u5_mult_82_CARRYB_15__31_,
         u5_mult_82_CARRYB_15__32_, u5_mult_82_CARRYB_15__33_,
         u5_mult_82_CARRYB_15__34_, u5_mult_82_CARRYB_15__35_,
         u5_mult_82_CARRYB_15__36_, u5_mult_82_CARRYB_15__37_,
         u5_mult_82_CARRYB_15__38_, u5_mult_82_CARRYB_15__39_,
         u5_mult_82_CARRYB_15__40_, u5_mult_82_CARRYB_15__41_,
         u5_mult_82_CARRYB_15__42_, u5_mult_82_CARRYB_15__43_,
         u5_mult_82_CARRYB_15__44_, u5_mult_82_CARRYB_15__45_,
         u5_mult_82_CARRYB_15__46_, u5_mult_82_CARRYB_15__47_,
         u5_mult_82_CARRYB_15__48_, u5_mult_82_CARRYB_15__49_,
         u5_mult_82_CARRYB_15__50_, u5_mult_82_CARRYB_15__51_,
         u5_mult_82_CARRYB_16__0_, u5_mult_82_CARRYB_16__1_,
         u5_mult_82_CARRYB_16__2_, u5_mult_82_CARRYB_16__3_,
         u5_mult_82_CARRYB_16__4_, u5_mult_82_CARRYB_16__5_,
         u5_mult_82_CARRYB_16__6_, u5_mult_82_CARRYB_16__7_,
         u5_mult_82_CARRYB_16__8_, u5_mult_82_CARRYB_16__9_,
         u5_mult_82_CARRYB_16__10_, u5_mult_82_CARRYB_16__11_,
         u5_mult_82_CARRYB_16__12_, u5_mult_82_CARRYB_16__13_,
         u5_mult_82_CARRYB_16__14_, u5_mult_82_CARRYB_16__15_,
         u5_mult_82_CARRYB_16__16_, u5_mult_82_CARRYB_16__17_,
         u5_mult_82_CARRYB_16__18_, u5_mult_82_CARRYB_16__19_,
         u5_mult_82_CARRYB_16__20_, u5_mult_82_CARRYB_16__21_,
         u5_mult_82_CARRYB_16__22_, u5_mult_82_CARRYB_16__23_,
         u5_mult_82_CARRYB_16__24_, u5_mult_82_CARRYB_16__25_,
         u5_mult_82_CARRYB_16__26_, u5_mult_82_CARRYB_16__27_,
         u5_mult_82_CARRYB_16__28_, u5_mult_82_CARRYB_16__29_,
         u5_mult_82_CARRYB_16__30_, u5_mult_82_CARRYB_16__31_,
         u5_mult_82_CARRYB_16__32_, u5_mult_82_CARRYB_16__33_,
         u5_mult_82_CARRYB_16__34_, u5_mult_82_CARRYB_16__35_,
         u5_mult_82_CARRYB_16__36_, u5_mult_82_CARRYB_16__37_,
         u5_mult_82_CARRYB_16__38_, u5_mult_82_CARRYB_16__39_,
         u5_mult_82_CARRYB_16__40_, u5_mult_82_CARRYB_16__41_,
         u5_mult_82_CARRYB_16__42_, u5_mult_82_CARRYB_16__43_,
         u5_mult_82_CARRYB_16__44_, u5_mult_82_CARRYB_16__45_,
         u5_mult_82_CARRYB_16__46_, u5_mult_82_CARRYB_16__47_,
         u5_mult_82_CARRYB_16__48_, u5_mult_82_CARRYB_16__49_,
         u5_mult_82_CARRYB_16__50_, u5_mult_82_CARRYB_16__51_,
         u5_mult_82_CARRYB_17__0_, u5_mult_82_CARRYB_17__1_,
         u5_mult_82_CARRYB_17__2_, u5_mult_82_CARRYB_17__3_,
         u5_mult_82_CARRYB_17__4_, u5_mult_82_CARRYB_17__5_,
         u5_mult_82_CARRYB_17__6_, u5_mult_82_CARRYB_17__7_,
         u5_mult_82_CARRYB_17__8_, u5_mult_82_CARRYB_17__9_,
         u5_mult_82_CARRYB_17__10_, u5_mult_82_CARRYB_17__11_,
         u5_mult_82_CARRYB_17__12_, u5_mult_82_CARRYB_17__13_,
         u5_mult_82_CARRYB_17__14_, u5_mult_82_CARRYB_17__15_,
         u5_mult_82_CARRYB_17__16_, u5_mult_82_CARRYB_17__17_,
         u5_mult_82_CARRYB_17__18_, u5_mult_82_CARRYB_17__19_,
         u5_mult_82_CARRYB_17__20_, u5_mult_82_CARRYB_17__21_,
         u5_mult_82_CARRYB_17__22_, u5_mult_82_CARRYB_17__23_,
         u5_mult_82_CARRYB_17__24_, u5_mult_82_CARRYB_17__25_,
         u5_mult_82_CARRYB_17__26_, u5_mult_82_CARRYB_17__27_,
         u5_mult_82_CARRYB_17__28_, u5_mult_82_CARRYB_17__29_,
         u5_mult_82_CARRYB_17__30_, u5_mult_82_CARRYB_17__31_,
         u5_mult_82_CARRYB_17__32_, u5_mult_82_CARRYB_17__33_,
         u5_mult_82_CARRYB_17__34_, u5_mult_82_CARRYB_17__35_,
         u5_mult_82_CARRYB_17__36_, u5_mult_82_CARRYB_17__37_,
         u5_mult_82_CARRYB_17__38_, u5_mult_82_CARRYB_17__39_,
         u5_mult_82_CARRYB_17__40_, u5_mult_82_CARRYB_17__41_,
         u5_mult_82_CARRYB_17__42_, u5_mult_82_CARRYB_17__43_,
         u5_mult_82_CARRYB_17__44_, u5_mult_82_CARRYB_17__45_,
         u5_mult_82_CARRYB_17__46_, u5_mult_82_CARRYB_17__47_,
         u5_mult_82_CARRYB_17__48_, u5_mult_82_CARRYB_17__49_,
         u5_mult_82_CARRYB_17__50_, u5_mult_82_CARRYB_17__51_,
         u5_mult_82_CARRYB_18__0_, u5_mult_82_CARRYB_18__1_,
         u5_mult_82_CARRYB_18__2_, u5_mult_82_CARRYB_18__3_,
         u5_mult_82_CARRYB_18__4_, u5_mult_82_CARRYB_18__5_,
         u5_mult_82_CARRYB_18__6_, u5_mult_82_CARRYB_18__7_,
         u5_mult_82_CARRYB_18__8_, u5_mult_82_CARRYB_18__9_,
         u5_mult_82_CARRYB_18__10_, u5_mult_82_CARRYB_18__11_,
         u5_mult_82_CARRYB_18__12_, u5_mult_82_CARRYB_18__13_,
         u5_mult_82_CARRYB_18__14_, u5_mult_82_CARRYB_18__15_,
         u5_mult_82_CARRYB_18__16_, u5_mult_82_CARRYB_18__17_,
         u5_mult_82_CARRYB_18__18_, u5_mult_82_CARRYB_18__19_,
         u5_mult_82_CARRYB_18__20_, u5_mult_82_CARRYB_18__21_,
         u5_mult_82_CARRYB_18__22_, u5_mult_82_CARRYB_18__23_,
         u5_mult_82_CARRYB_18__24_, u5_mult_82_CARRYB_18__25_,
         u5_mult_82_CARRYB_18__26_, u5_mult_82_CARRYB_18__27_,
         u5_mult_82_CARRYB_18__28_, u5_mult_82_CARRYB_18__29_,
         u5_mult_82_CARRYB_18__30_, u5_mult_82_CARRYB_18__31_,
         u5_mult_82_CARRYB_18__32_, u5_mult_82_CARRYB_18__33_,
         u5_mult_82_CARRYB_18__34_, u5_mult_82_CARRYB_18__35_,
         u5_mult_82_CARRYB_18__36_, u5_mult_82_CARRYB_18__37_,
         u5_mult_82_CARRYB_18__38_, u5_mult_82_CARRYB_18__39_,
         u5_mult_82_CARRYB_18__40_, u5_mult_82_CARRYB_18__41_,
         u5_mult_82_CARRYB_18__42_, u5_mult_82_CARRYB_18__43_,
         u5_mult_82_CARRYB_18__44_, u5_mult_82_CARRYB_18__45_,
         u5_mult_82_CARRYB_18__46_, u5_mult_82_CARRYB_18__47_,
         u5_mult_82_CARRYB_18__48_, u5_mult_82_CARRYB_18__49_,
         u5_mult_82_CARRYB_18__50_, u5_mult_82_CARRYB_18__51_,
         u5_mult_82_CARRYB_19__0_, u5_mult_82_CARRYB_19__1_,
         u5_mult_82_CARRYB_19__2_, u5_mult_82_CARRYB_19__3_,
         u5_mult_82_CARRYB_19__4_, u5_mult_82_CARRYB_19__5_,
         u5_mult_82_CARRYB_19__6_, u5_mult_82_CARRYB_19__7_,
         u5_mult_82_CARRYB_19__8_, u5_mult_82_CARRYB_19__9_,
         u5_mult_82_CARRYB_19__10_, u5_mult_82_CARRYB_19__11_,
         u5_mult_82_CARRYB_19__12_, u5_mult_82_CARRYB_19__13_,
         u5_mult_82_CARRYB_19__14_, u5_mult_82_CARRYB_19__15_,
         u5_mult_82_CARRYB_19__16_, u5_mult_82_CARRYB_19__17_,
         u5_mult_82_CARRYB_19__18_, u5_mult_82_CARRYB_19__19_,
         u5_mult_82_CARRYB_19__20_, u5_mult_82_CARRYB_19__21_,
         u5_mult_82_CARRYB_19__22_, u5_mult_82_CARRYB_19__23_,
         u5_mult_82_CARRYB_19__24_, u5_mult_82_CARRYB_19__25_,
         u5_mult_82_CARRYB_19__26_, u5_mult_82_CARRYB_19__27_,
         u5_mult_82_CARRYB_19__28_, u5_mult_82_CARRYB_19__29_,
         u5_mult_82_CARRYB_19__30_, u5_mult_82_CARRYB_19__31_,
         u5_mult_82_CARRYB_19__32_, u5_mult_82_CARRYB_19__33_,
         u5_mult_82_CARRYB_19__34_, u5_mult_82_CARRYB_19__35_,
         u5_mult_82_CARRYB_19__36_, u5_mult_82_CARRYB_19__37_,
         u5_mult_82_CARRYB_19__38_, u5_mult_82_CARRYB_19__39_,
         u5_mult_82_CARRYB_19__40_, u5_mult_82_CARRYB_19__41_,
         u5_mult_82_CARRYB_19__42_, u5_mult_82_CARRYB_19__43_,
         u5_mult_82_CARRYB_19__44_, u5_mult_82_CARRYB_19__45_,
         u5_mult_82_CARRYB_19__46_, u5_mult_82_CARRYB_19__47_,
         u5_mult_82_CARRYB_19__48_, u5_mult_82_CARRYB_19__49_,
         u5_mult_82_CARRYB_19__50_, u5_mult_82_CARRYB_19__51_,
         u5_mult_82_CARRYB_20__0_, u5_mult_82_CARRYB_20__1_,
         u5_mult_82_CARRYB_20__2_, u5_mult_82_CARRYB_20__3_,
         u5_mult_82_CARRYB_20__4_, u5_mult_82_CARRYB_20__5_,
         u5_mult_82_CARRYB_20__6_, u5_mult_82_CARRYB_20__7_,
         u5_mult_82_CARRYB_20__8_, u5_mult_82_CARRYB_20__9_,
         u5_mult_82_CARRYB_20__10_, u5_mult_82_CARRYB_20__11_,
         u5_mult_82_CARRYB_20__12_, u5_mult_82_CARRYB_20__13_,
         u5_mult_82_CARRYB_20__14_, u5_mult_82_CARRYB_20__15_,
         u5_mult_82_CARRYB_20__16_, u5_mult_82_CARRYB_20__17_,
         u5_mult_82_CARRYB_20__18_, u5_mult_82_CARRYB_20__19_,
         u5_mult_82_CARRYB_20__20_, u5_mult_82_CARRYB_20__21_,
         u5_mult_82_CARRYB_20__22_, u5_mult_82_CARRYB_20__23_,
         u5_mult_82_CARRYB_20__24_, u5_mult_82_CARRYB_20__25_,
         u5_mult_82_CARRYB_20__26_, u5_mult_82_CARRYB_20__27_,
         u5_mult_82_CARRYB_20__28_, u5_mult_82_CARRYB_20__29_,
         u5_mult_82_CARRYB_20__30_, u5_mult_82_CARRYB_20__31_,
         u5_mult_82_CARRYB_20__32_, u5_mult_82_CARRYB_20__33_,
         u5_mult_82_CARRYB_20__34_, u5_mult_82_CARRYB_20__35_,
         u5_mult_82_CARRYB_20__36_, u5_mult_82_CARRYB_20__37_,
         u5_mult_82_CARRYB_20__38_, u5_mult_82_CARRYB_20__39_,
         u5_mult_82_CARRYB_20__40_, u5_mult_82_CARRYB_20__41_,
         u5_mult_82_CARRYB_20__42_, u5_mult_82_CARRYB_20__43_,
         u5_mult_82_CARRYB_20__44_, u5_mult_82_CARRYB_20__45_,
         u5_mult_82_CARRYB_20__46_, u5_mult_82_CARRYB_20__47_,
         u5_mult_82_CARRYB_20__48_, u5_mult_82_CARRYB_20__49_,
         u5_mult_82_CARRYB_20__50_, u5_mult_82_CARRYB_20__51_,
         u5_mult_82_CARRYB_21__0_, u5_mult_82_CARRYB_21__1_,
         u5_mult_82_CARRYB_21__2_, u5_mult_82_CARRYB_21__3_,
         u5_mult_82_CARRYB_21__4_, u5_mult_82_CARRYB_21__5_,
         u5_mult_82_CARRYB_21__6_, u5_mult_82_CARRYB_21__7_,
         u5_mult_82_CARRYB_21__8_, u5_mult_82_CARRYB_21__9_,
         u5_mult_82_CARRYB_21__10_, u5_mult_82_CARRYB_21__11_,
         u5_mult_82_CARRYB_21__12_, u5_mult_82_CARRYB_21__13_,
         u5_mult_82_CARRYB_21__14_, u5_mult_82_CARRYB_21__15_,
         u5_mult_82_CARRYB_21__16_, u5_mult_82_CARRYB_21__17_,
         u5_mult_82_CARRYB_21__18_, u5_mult_82_CARRYB_21__19_,
         u5_mult_82_CARRYB_21__20_, u5_mult_82_CARRYB_21__21_,
         u5_mult_82_CARRYB_21__22_, u5_mult_82_CARRYB_21__23_,
         u5_mult_82_CARRYB_21__24_, u5_mult_82_CARRYB_21__25_,
         u5_mult_82_CARRYB_21__26_, u5_mult_82_CARRYB_21__27_,
         u5_mult_82_CARRYB_21__28_, u5_mult_82_CARRYB_21__29_,
         u5_mult_82_CARRYB_21__30_, u5_mult_82_CARRYB_21__31_,
         u5_mult_82_CARRYB_21__32_, u5_mult_82_CARRYB_21__33_,
         u5_mult_82_CARRYB_21__34_, u5_mult_82_CARRYB_21__35_,
         u5_mult_82_CARRYB_21__36_, u5_mult_82_CARRYB_21__37_,
         u5_mult_82_CARRYB_21__38_, u5_mult_82_CARRYB_21__39_,
         u5_mult_82_CARRYB_21__40_, u5_mult_82_CARRYB_21__41_,
         u5_mult_82_CARRYB_21__42_, u5_mult_82_CARRYB_21__43_,
         u5_mult_82_CARRYB_21__44_, u5_mult_82_CARRYB_21__45_,
         u5_mult_82_CARRYB_21__46_, u5_mult_82_CARRYB_21__47_,
         u5_mult_82_CARRYB_21__48_, u5_mult_82_CARRYB_21__49_,
         u5_mult_82_CARRYB_21__50_, u5_mult_82_CARRYB_21__51_,
         u5_mult_82_CARRYB_22__0_, u5_mult_82_CARRYB_22__1_,
         u5_mult_82_CARRYB_22__2_, u5_mult_82_CARRYB_22__3_,
         u5_mult_82_CARRYB_22__4_, u5_mult_82_CARRYB_22__5_,
         u5_mult_82_CARRYB_22__6_, u5_mult_82_CARRYB_22__7_,
         u5_mult_82_CARRYB_22__8_, u5_mult_82_CARRYB_22__9_,
         u5_mult_82_CARRYB_22__10_, u5_mult_82_CARRYB_22__11_,
         u5_mult_82_CARRYB_22__12_, u5_mult_82_CARRYB_22__13_,
         u5_mult_82_CARRYB_22__14_, u5_mult_82_CARRYB_22__15_,
         u5_mult_82_CARRYB_22__16_, u5_mult_82_CARRYB_22__17_,
         u5_mult_82_CARRYB_22__18_, u5_mult_82_CARRYB_22__19_,
         u5_mult_82_CARRYB_22__20_, u5_mult_82_CARRYB_22__21_,
         u5_mult_82_CARRYB_22__22_, u5_mult_82_CARRYB_22__23_,
         u5_mult_82_CARRYB_22__24_, u5_mult_82_CARRYB_22__25_,
         u5_mult_82_CARRYB_22__26_, u5_mult_82_CARRYB_22__27_,
         u5_mult_82_CARRYB_22__28_, u5_mult_82_CARRYB_22__29_,
         u5_mult_82_CARRYB_22__30_, u5_mult_82_CARRYB_22__31_,
         u5_mult_82_CARRYB_22__32_, u5_mult_82_CARRYB_22__33_,
         u5_mult_82_CARRYB_22__34_, u5_mult_82_CARRYB_22__35_,
         u5_mult_82_CARRYB_22__36_, u5_mult_82_CARRYB_22__37_,
         u5_mult_82_CARRYB_22__38_, u5_mult_82_CARRYB_22__39_,
         u5_mult_82_CARRYB_22__40_, u5_mult_82_CARRYB_22__41_,
         u5_mult_82_CARRYB_22__42_, u5_mult_82_CARRYB_22__43_,
         u5_mult_82_CARRYB_22__44_, u5_mult_82_CARRYB_22__45_,
         u5_mult_82_CARRYB_22__46_, u5_mult_82_CARRYB_22__47_,
         u5_mult_82_CARRYB_22__48_, u5_mult_82_CARRYB_22__49_,
         u5_mult_82_CARRYB_22__50_, u5_mult_82_CARRYB_22__51_,
         u5_mult_82_CARRYB_23__0_, u5_mult_82_CARRYB_23__1_,
         u5_mult_82_CARRYB_23__2_, u5_mult_82_CARRYB_23__3_,
         u5_mult_82_CARRYB_23__4_, u5_mult_82_CARRYB_23__5_,
         u5_mult_82_CARRYB_23__6_, u5_mult_82_CARRYB_23__7_,
         u5_mult_82_CARRYB_23__8_, u5_mult_82_CARRYB_23__9_,
         u5_mult_82_CARRYB_23__10_, u5_mult_82_CARRYB_23__11_,
         u5_mult_82_CARRYB_23__12_, u5_mult_82_CARRYB_23__13_,
         u5_mult_82_CARRYB_23__14_, u5_mult_82_CARRYB_23__15_,
         u5_mult_82_CARRYB_23__16_, u5_mult_82_CARRYB_23__17_,
         u5_mult_82_CARRYB_23__18_, u5_mult_82_CARRYB_23__19_,
         u5_mult_82_CARRYB_23__20_, u5_mult_82_CARRYB_23__21_,
         u5_mult_82_CARRYB_23__22_, u5_mult_82_CARRYB_23__23_,
         u5_mult_82_CARRYB_23__24_, u5_mult_82_CARRYB_23__25_,
         u5_mult_82_CARRYB_23__26_, u5_mult_82_CARRYB_23__27_,
         u5_mult_82_CARRYB_23__28_, u5_mult_82_CARRYB_23__29_,
         u5_mult_82_CARRYB_23__30_, u5_mult_82_CARRYB_23__31_,
         u5_mult_82_CARRYB_23__32_, u5_mult_82_CARRYB_23__33_,
         u5_mult_82_CARRYB_23__34_, u5_mult_82_CARRYB_23__35_,
         u5_mult_82_CARRYB_23__36_, u5_mult_82_CARRYB_23__37_,
         u5_mult_82_CARRYB_23__38_, u5_mult_82_CARRYB_23__39_,
         u5_mult_82_CARRYB_23__40_, u5_mult_82_CARRYB_23__41_,
         u5_mult_82_CARRYB_23__42_, u5_mult_82_CARRYB_23__43_,
         u5_mult_82_CARRYB_23__44_, u5_mult_82_CARRYB_23__45_,
         u5_mult_82_CARRYB_23__46_, u5_mult_82_CARRYB_23__47_,
         u5_mult_82_CARRYB_23__48_, u5_mult_82_CARRYB_23__49_,
         u5_mult_82_CARRYB_23__50_, u5_mult_82_CARRYB_23__51_,
         u5_mult_82_CARRYB_24__0_, u5_mult_82_SUMB_4__37_,
         u5_mult_82_SUMB_4__38_, u5_mult_82_SUMB_4__39_,
         u5_mult_82_SUMB_4__40_, u5_mult_82_SUMB_4__41_,
         u5_mult_82_SUMB_4__42_, u5_mult_82_SUMB_4__43_,
         u5_mult_82_SUMB_4__44_, u5_mult_82_SUMB_4__45_,
         u5_mult_82_SUMB_4__46_, u5_mult_82_SUMB_4__47_,
         u5_mult_82_SUMB_4__48_, u5_mult_82_SUMB_4__49_,
         u5_mult_82_SUMB_4__50_, u5_mult_82_SUMB_4__51_, u5_mult_82_SUMB_5__1_,
         u5_mult_82_SUMB_5__2_, u5_mult_82_SUMB_5__3_, u5_mult_82_SUMB_5__4_,
         u5_mult_82_SUMB_5__5_, u5_mult_82_SUMB_5__6_, u5_mult_82_SUMB_5__7_,
         u5_mult_82_SUMB_5__8_, u5_mult_82_SUMB_5__9_, u5_mult_82_SUMB_5__10_,
         u5_mult_82_SUMB_5__11_, u5_mult_82_SUMB_5__12_,
         u5_mult_82_SUMB_5__13_, u5_mult_82_SUMB_5__14_,
         u5_mult_82_SUMB_5__15_, u5_mult_82_SUMB_5__16_,
         u5_mult_82_SUMB_5__17_, u5_mult_82_SUMB_5__18_,
         u5_mult_82_SUMB_5__19_, u5_mult_82_SUMB_5__20_,
         u5_mult_82_SUMB_5__21_, u5_mult_82_SUMB_5__22_,
         u5_mult_82_SUMB_5__23_, u5_mult_82_SUMB_5__24_,
         u5_mult_82_SUMB_5__25_, u5_mult_82_SUMB_5__26_,
         u5_mult_82_SUMB_5__27_, u5_mult_82_SUMB_5__28_,
         u5_mult_82_SUMB_5__29_, u5_mult_82_SUMB_5__30_,
         u5_mult_82_SUMB_5__31_, u5_mult_82_SUMB_5__32_,
         u5_mult_82_SUMB_5__33_, u5_mult_82_SUMB_5__34_,
         u5_mult_82_SUMB_5__35_, u5_mult_82_SUMB_5__36_,
         u5_mult_82_SUMB_5__37_, u5_mult_82_SUMB_5__38_,
         u5_mult_82_SUMB_5__39_, u5_mult_82_SUMB_5__40_,
         u5_mult_82_SUMB_5__41_, u5_mult_82_SUMB_5__42_,
         u5_mult_82_SUMB_5__43_, u5_mult_82_SUMB_5__44_,
         u5_mult_82_SUMB_5__45_, u5_mult_82_SUMB_5__46_,
         u5_mult_82_SUMB_5__47_, u5_mult_82_SUMB_5__48_,
         u5_mult_82_SUMB_5__49_, u5_mult_82_SUMB_5__50_,
         u5_mult_82_SUMB_5__51_, u5_mult_82_SUMB_6__1_, u5_mult_82_SUMB_6__2_,
         u5_mult_82_SUMB_6__3_, u5_mult_82_SUMB_6__4_, u5_mult_82_SUMB_6__5_,
         u5_mult_82_SUMB_6__6_, u5_mult_82_SUMB_6__7_, u5_mult_82_SUMB_6__8_,
         u5_mult_82_SUMB_6__9_, u5_mult_82_SUMB_6__10_, u5_mult_82_SUMB_6__11_,
         u5_mult_82_SUMB_6__12_, u5_mult_82_SUMB_6__13_,
         u5_mult_82_SUMB_6__14_, u5_mult_82_SUMB_6__15_,
         u5_mult_82_SUMB_6__16_, u5_mult_82_SUMB_6__17_,
         u5_mult_82_SUMB_6__18_, u5_mult_82_SUMB_6__19_,
         u5_mult_82_SUMB_6__20_, u5_mult_82_SUMB_6__21_,
         u5_mult_82_SUMB_6__22_, u5_mult_82_SUMB_6__23_,
         u5_mult_82_SUMB_6__24_, u5_mult_82_SUMB_6__25_,
         u5_mult_82_SUMB_6__26_, u5_mult_82_SUMB_6__27_,
         u5_mult_82_SUMB_6__28_, u5_mult_82_SUMB_6__29_,
         u5_mult_82_SUMB_6__30_, u5_mult_82_SUMB_6__31_,
         u5_mult_82_SUMB_6__32_, u5_mult_82_SUMB_6__33_,
         u5_mult_82_SUMB_6__34_, u5_mult_82_SUMB_6__35_,
         u5_mult_82_SUMB_6__36_, u5_mult_82_SUMB_6__37_,
         u5_mult_82_SUMB_6__38_, u5_mult_82_SUMB_6__39_,
         u5_mult_82_SUMB_6__40_, u5_mult_82_SUMB_6__41_,
         u5_mult_82_SUMB_6__42_, u5_mult_82_SUMB_6__43_,
         u5_mult_82_SUMB_6__44_, u5_mult_82_SUMB_6__45_,
         u5_mult_82_SUMB_6__46_, u5_mult_82_SUMB_6__47_,
         u5_mult_82_SUMB_6__48_, u5_mult_82_SUMB_6__49_,
         u5_mult_82_SUMB_6__50_, u5_mult_82_SUMB_6__51_, u5_mult_82_SUMB_7__1_,
         u5_mult_82_SUMB_7__2_, u5_mult_82_SUMB_7__3_, u5_mult_82_SUMB_7__4_,
         u5_mult_82_SUMB_7__5_, u5_mult_82_SUMB_7__6_, u5_mult_82_SUMB_7__7_,
         u5_mult_82_SUMB_7__8_, u5_mult_82_SUMB_7__9_, u5_mult_82_SUMB_7__10_,
         u5_mult_82_SUMB_7__11_, u5_mult_82_SUMB_7__12_,
         u5_mult_82_SUMB_7__13_, u5_mult_82_SUMB_7__14_,
         u5_mult_82_SUMB_7__15_, u5_mult_82_SUMB_7__16_,
         u5_mult_82_SUMB_7__17_, u5_mult_82_SUMB_7__18_,
         u5_mult_82_SUMB_7__19_, u5_mult_82_SUMB_7__20_,
         u5_mult_82_SUMB_7__21_, u5_mult_82_SUMB_7__22_,
         u5_mult_82_SUMB_7__23_, u5_mult_82_SUMB_7__24_,
         u5_mult_82_SUMB_7__25_, u5_mult_82_SUMB_7__26_,
         u5_mult_82_SUMB_7__27_, u5_mult_82_SUMB_7__28_,
         u5_mult_82_SUMB_7__29_, u5_mult_82_SUMB_7__30_,
         u5_mult_82_SUMB_7__31_, u5_mult_82_SUMB_7__32_,
         u5_mult_82_SUMB_7__33_, u5_mult_82_SUMB_7__34_,
         u5_mult_82_SUMB_7__35_, u5_mult_82_SUMB_7__36_,
         u5_mult_82_SUMB_7__37_, u5_mult_82_SUMB_7__38_,
         u5_mult_82_SUMB_7__39_, u5_mult_82_SUMB_7__40_,
         u5_mult_82_SUMB_7__41_, u5_mult_82_SUMB_7__42_,
         u5_mult_82_SUMB_7__43_, u5_mult_82_SUMB_7__44_,
         u5_mult_82_SUMB_7__45_, u5_mult_82_SUMB_7__46_,
         u5_mult_82_SUMB_7__47_, u5_mult_82_SUMB_7__48_,
         u5_mult_82_SUMB_7__49_, u5_mult_82_SUMB_7__50_,
         u5_mult_82_SUMB_7__51_, u5_mult_82_SUMB_8__1_, u5_mult_82_SUMB_8__2_,
         u5_mult_82_SUMB_8__3_, u5_mult_82_SUMB_8__4_, u5_mult_82_SUMB_8__5_,
         u5_mult_82_SUMB_8__6_, u5_mult_82_SUMB_8__7_, u5_mult_82_SUMB_8__8_,
         u5_mult_82_SUMB_8__9_, u5_mult_82_SUMB_8__10_, u5_mult_82_SUMB_8__11_,
         u5_mult_82_SUMB_8__12_, u5_mult_82_SUMB_8__13_,
         u5_mult_82_SUMB_8__14_, u5_mult_82_SUMB_8__15_,
         u5_mult_82_SUMB_8__16_, u5_mult_82_SUMB_8__17_,
         u5_mult_82_SUMB_8__18_, u5_mult_82_SUMB_8__19_,
         u5_mult_82_SUMB_8__20_, u5_mult_82_SUMB_8__21_,
         u5_mult_82_SUMB_8__22_, u5_mult_82_SUMB_8__23_,
         u5_mult_82_SUMB_8__24_, u5_mult_82_SUMB_8__25_,
         u5_mult_82_SUMB_8__26_, u5_mult_82_SUMB_8__27_,
         u5_mult_82_SUMB_8__28_, u5_mult_82_SUMB_8__29_,
         u5_mult_82_SUMB_8__30_, u5_mult_82_SUMB_8__31_,
         u5_mult_82_SUMB_8__32_, u5_mult_82_SUMB_8__33_,
         u5_mult_82_SUMB_8__34_, u5_mult_82_SUMB_8__35_,
         u5_mult_82_SUMB_8__36_, u5_mult_82_SUMB_8__37_,
         u5_mult_82_SUMB_8__38_, u5_mult_82_SUMB_8__39_,
         u5_mult_82_SUMB_8__40_, u5_mult_82_SUMB_8__41_,
         u5_mult_82_SUMB_8__42_, u5_mult_82_SUMB_8__43_,
         u5_mult_82_SUMB_8__44_, u5_mult_82_SUMB_8__45_,
         u5_mult_82_SUMB_8__46_, u5_mult_82_SUMB_8__47_,
         u5_mult_82_SUMB_8__48_, u5_mult_82_SUMB_8__49_,
         u5_mult_82_SUMB_8__50_, u5_mult_82_SUMB_8__51_, u5_mult_82_SUMB_9__1_,
         u5_mult_82_SUMB_9__2_, u5_mult_82_SUMB_9__3_, u5_mult_82_SUMB_9__4_,
         u5_mult_82_SUMB_9__5_, u5_mult_82_SUMB_9__6_, u5_mult_82_SUMB_9__7_,
         u5_mult_82_SUMB_9__8_, u5_mult_82_SUMB_9__9_, u5_mult_82_SUMB_9__10_,
         u5_mult_82_SUMB_9__11_, u5_mult_82_SUMB_9__12_,
         u5_mult_82_SUMB_9__13_, u5_mult_82_SUMB_9__14_,
         u5_mult_82_SUMB_9__15_, u5_mult_82_SUMB_9__16_,
         u5_mult_82_SUMB_9__17_, u5_mult_82_SUMB_9__18_,
         u5_mult_82_SUMB_9__19_, u5_mult_82_SUMB_9__20_,
         u5_mult_82_SUMB_9__21_, u5_mult_82_SUMB_9__22_,
         u5_mult_82_SUMB_9__23_, u5_mult_82_SUMB_9__24_,
         u5_mult_82_SUMB_9__25_, u5_mult_82_SUMB_9__26_,
         u5_mult_82_SUMB_9__27_, u5_mult_82_SUMB_9__28_,
         u5_mult_82_SUMB_9__29_, u5_mult_82_SUMB_9__30_,
         u5_mult_82_SUMB_9__31_, u5_mult_82_SUMB_9__32_,
         u5_mult_82_SUMB_9__33_, u5_mult_82_SUMB_9__34_,
         u5_mult_82_SUMB_9__35_, u5_mult_82_SUMB_9__36_,
         u5_mult_82_SUMB_9__37_, u5_mult_82_SUMB_9__38_,
         u5_mult_82_SUMB_9__39_, u5_mult_82_SUMB_9__40_,
         u5_mult_82_SUMB_9__41_, u5_mult_82_SUMB_9__42_,
         u5_mult_82_SUMB_9__43_, u5_mult_82_SUMB_9__44_,
         u5_mult_82_SUMB_9__45_, u5_mult_82_SUMB_9__46_,
         u5_mult_82_SUMB_9__47_, u5_mult_82_SUMB_9__48_,
         u5_mult_82_SUMB_9__49_, u5_mult_82_SUMB_9__50_,
         u5_mult_82_SUMB_9__51_, u5_mult_82_SUMB_10__1_,
         u5_mult_82_SUMB_10__2_, u5_mult_82_SUMB_10__3_,
         u5_mult_82_SUMB_10__4_, u5_mult_82_SUMB_10__5_,
         u5_mult_82_SUMB_10__6_, u5_mult_82_SUMB_10__7_,
         u5_mult_82_SUMB_10__8_, u5_mult_82_SUMB_10__9_,
         u5_mult_82_SUMB_10__10_, u5_mult_82_SUMB_10__11_,
         u5_mult_82_SUMB_10__12_, u5_mult_82_SUMB_10__13_,
         u5_mult_82_SUMB_10__14_, u5_mult_82_SUMB_10__15_,
         u5_mult_82_SUMB_10__16_, u5_mult_82_SUMB_10__17_,
         u5_mult_82_SUMB_10__18_, u5_mult_82_SUMB_10__19_,
         u5_mult_82_SUMB_10__20_, u5_mult_82_SUMB_10__21_,
         u5_mult_82_SUMB_10__22_, u5_mult_82_SUMB_10__23_,
         u5_mult_82_SUMB_10__24_, u5_mult_82_SUMB_10__25_,
         u5_mult_82_SUMB_10__26_, u5_mult_82_SUMB_10__27_,
         u5_mult_82_SUMB_10__28_, u5_mult_82_SUMB_10__29_,
         u5_mult_82_SUMB_10__30_, u5_mult_82_SUMB_10__31_,
         u5_mult_82_SUMB_10__32_, u5_mult_82_SUMB_10__33_,
         u5_mult_82_SUMB_10__34_, u5_mult_82_SUMB_10__35_,
         u5_mult_82_SUMB_10__36_, u5_mult_82_SUMB_10__37_,
         u5_mult_82_SUMB_10__38_, u5_mult_82_SUMB_10__39_,
         u5_mult_82_SUMB_10__40_, u5_mult_82_SUMB_10__41_,
         u5_mult_82_SUMB_10__42_, u5_mult_82_SUMB_10__43_,
         u5_mult_82_SUMB_10__44_, u5_mult_82_SUMB_10__45_,
         u5_mult_82_SUMB_10__46_, u5_mult_82_SUMB_10__47_,
         u5_mult_82_SUMB_10__48_, u5_mult_82_SUMB_10__49_,
         u5_mult_82_SUMB_10__50_, u5_mult_82_SUMB_10__51_,
         u5_mult_82_SUMB_11__1_, u5_mult_82_SUMB_11__2_,
         u5_mult_82_SUMB_11__3_, u5_mult_82_SUMB_11__4_,
         u5_mult_82_SUMB_11__5_, u5_mult_82_SUMB_11__6_,
         u5_mult_82_SUMB_11__7_, u5_mult_82_SUMB_11__8_,
         u5_mult_82_SUMB_11__9_, u5_mult_82_SUMB_11__10_,
         u5_mult_82_SUMB_11__11_, u5_mult_82_SUMB_11__12_,
         u5_mult_82_SUMB_11__13_, u5_mult_82_SUMB_11__14_,
         u5_mult_82_SUMB_11__15_, u5_mult_82_SUMB_11__16_,
         u5_mult_82_SUMB_11__17_, u5_mult_82_SUMB_11__18_,
         u5_mult_82_SUMB_11__19_, u5_mult_82_SUMB_11__20_,
         u5_mult_82_SUMB_11__21_, u5_mult_82_SUMB_11__22_,
         u5_mult_82_SUMB_11__23_, u5_mult_82_SUMB_11__24_,
         u5_mult_82_SUMB_11__25_, u5_mult_82_SUMB_11__26_,
         u5_mult_82_SUMB_11__27_, u5_mult_82_SUMB_11__28_,
         u5_mult_82_SUMB_11__29_, u5_mult_82_SUMB_11__30_,
         u5_mult_82_SUMB_11__31_, u5_mult_82_SUMB_11__32_,
         u5_mult_82_SUMB_11__33_, u5_mult_82_SUMB_11__34_,
         u5_mult_82_SUMB_11__35_, u5_mult_82_SUMB_11__36_,
         u5_mult_82_SUMB_11__37_, u5_mult_82_SUMB_11__38_,
         u5_mult_82_SUMB_11__39_, u5_mult_82_SUMB_11__40_,
         u5_mult_82_SUMB_11__41_, u5_mult_82_SUMB_11__42_,
         u5_mult_82_SUMB_11__43_, u5_mult_82_SUMB_11__44_,
         u5_mult_82_SUMB_11__45_, u5_mult_82_SUMB_11__46_,
         u5_mult_82_SUMB_11__47_, u5_mult_82_SUMB_11__48_,
         u5_mult_82_SUMB_11__49_, u5_mult_82_SUMB_11__50_,
         u5_mult_82_SUMB_11__51_, u5_mult_82_SUMB_12__1_,
         u5_mult_82_SUMB_12__2_, u5_mult_82_SUMB_12__3_,
         u5_mult_82_SUMB_12__4_, u5_mult_82_SUMB_12__5_,
         u5_mult_82_SUMB_12__6_, u5_mult_82_SUMB_12__7_,
         u5_mult_82_SUMB_12__8_, u5_mult_82_SUMB_12__9_,
         u5_mult_82_SUMB_12__10_, u5_mult_82_SUMB_12__11_,
         u5_mult_82_SUMB_12__12_, u5_mult_82_SUMB_12__13_,
         u5_mult_82_SUMB_12__14_, u5_mult_82_SUMB_12__15_,
         u5_mult_82_SUMB_12__16_, u5_mult_82_SUMB_12__17_,
         u5_mult_82_SUMB_12__18_, u5_mult_82_SUMB_12__19_,
         u5_mult_82_SUMB_12__20_, u5_mult_82_SUMB_12__21_,
         u5_mult_82_SUMB_12__22_, u5_mult_82_SUMB_12__23_,
         u5_mult_82_SUMB_12__24_, u5_mult_82_SUMB_12__25_,
         u5_mult_82_SUMB_12__26_, u5_mult_82_SUMB_12__27_,
         u5_mult_82_SUMB_12__28_, u5_mult_82_SUMB_12__29_,
         u5_mult_82_SUMB_12__30_, u5_mult_82_SUMB_12__31_,
         u5_mult_82_SUMB_12__32_, u5_mult_82_SUMB_12__33_,
         u5_mult_82_SUMB_12__34_, u5_mult_82_SUMB_12__35_,
         u5_mult_82_SUMB_12__36_, u5_mult_82_SUMB_12__37_,
         u5_mult_82_SUMB_12__38_, u5_mult_82_SUMB_12__39_,
         u5_mult_82_SUMB_12__40_, u5_mult_82_SUMB_12__41_,
         u5_mult_82_SUMB_12__42_, u5_mult_82_SUMB_12__43_,
         u5_mult_82_SUMB_12__44_, u5_mult_82_SUMB_12__45_,
         u5_mult_82_SUMB_12__46_, u5_mult_82_SUMB_12__47_,
         u5_mult_82_SUMB_12__48_, u5_mult_82_SUMB_12__49_,
         u5_mult_82_SUMB_12__50_, u5_mult_82_SUMB_12__51_,
         u5_mult_82_SUMB_13__1_, u5_mult_82_SUMB_13__2_,
         u5_mult_82_SUMB_13__3_, u5_mult_82_SUMB_13__4_,
         u5_mult_82_SUMB_13__5_, u5_mult_82_SUMB_13__6_,
         u5_mult_82_SUMB_13__7_, u5_mult_82_SUMB_13__8_,
         u5_mult_82_SUMB_13__9_, u5_mult_82_SUMB_13__10_,
         u5_mult_82_SUMB_13__11_, u5_mult_82_SUMB_13__12_,
         u5_mult_82_SUMB_13__13_, u5_mult_82_SUMB_13__14_,
         u5_mult_82_SUMB_13__15_, u5_mult_82_SUMB_13__16_,
         u5_mult_82_SUMB_13__17_, u5_mult_82_SUMB_13__18_,
         u5_mult_82_SUMB_13__19_, u5_mult_82_SUMB_13__20_,
         u5_mult_82_SUMB_13__21_, u5_mult_82_SUMB_13__22_,
         u5_mult_82_SUMB_13__23_, u5_mult_82_SUMB_13__24_,
         u5_mult_82_SUMB_13__25_, u5_mult_82_SUMB_13__26_,
         u5_mult_82_SUMB_13__27_, u5_mult_82_SUMB_13__28_,
         u5_mult_82_SUMB_13__29_, u5_mult_82_SUMB_13__30_,
         u5_mult_82_SUMB_13__31_, u5_mult_82_SUMB_13__32_,
         u5_mult_82_SUMB_13__33_, u5_mult_82_SUMB_13__34_,
         u5_mult_82_SUMB_13__35_, u5_mult_82_SUMB_13__36_,
         u5_mult_82_SUMB_13__37_, u5_mult_82_SUMB_13__38_,
         u5_mult_82_SUMB_13__39_, u5_mult_82_SUMB_13__40_,
         u5_mult_82_SUMB_13__41_, u5_mult_82_SUMB_13__42_,
         u5_mult_82_SUMB_13__43_, u5_mult_82_SUMB_13__44_,
         u5_mult_82_SUMB_13__45_, u5_mult_82_SUMB_13__46_,
         u5_mult_82_SUMB_13__47_, u5_mult_82_SUMB_13__48_,
         u5_mult_82_SUMB_13__49_, u5_mult_82_SUMB_13__50_,
         u5_mult_82_SUMB_13__51_, u5_mult_82_SUMB_14__1_,
         u5_mult_82_SUMB_14__2_, u5_mult_82_SUMB_14__3_,
         u5_mult_82_SUMB_14__4_, u5_mult_82_SUMB_14__5_,
         u5_mult_82_SUMB_14__6_, u5_mult_82_SUMB_14__7_,
         u5_mult_82_SUMB_14__8_, u5_mult_82_SUMB_14__9_,
         u5_mult_82_SUMB_14__10_, u5_mult_82_SUMB_14__11_,
         u5_mult_82_SUMB_14__12_, u5_mult_82_SUMB_14__13_,
         u5_mult_82_SUMB_14__14_, u5_mult_82_SUMB_14__15_,
         u5_mult_82_SUMB_14__16_, u5_mult_82_SUMB_14__17_,
         u5_mult_82_SUMB_14__18_, u5_mult_82_CARRYB_4__37_,
         u5_mult_82_CARRYB_4__38_, u5_mult_82_CARRYB_4__39_,
         u5_mult_82_CARRYB_4__40_, u5_mult_82_CARRYB_4__41_,
         u5_mult_82_CARRYB_4__42_, u5_mult_82_CARRYB_4__43_,
         u5_mult_82_CARRYB_4__44_, u5_mult_82_CARRYB_4__45_,
         u5_mult_82_CARRYB_4__46_, u5_mult_82_CARRYB_4__47_,
         u5_mult_82_CARRYB_4__48_, u5_mult_82_CARRYB_4__49_,
         u5_mult_82_CARRYB_4__50_, u5_mult_82_CARRYB_4__51_,
         u5_mult_82_CARRYB_5__0_, u5_mult_82_CARRYB_5__1_,
         u5_mult_82_CARRYB_5__2_, u5_mult_82_CARRYB_5__3_,
         u5_mult_82_CARRYB_5__4_, u5_mult_82_CARRYB_5__5_,
         u5_mult_82_CARRYB_5__6_, u5_mult_82_CARRYB_5__7_,
         u5_mult_82_CARRYB_5__8_, u5_mult_82_CARRYB_5__9_,
         u5_mult_82_CARRYB_5__10_, u5_mult_82_CARRYB_5__11_,
         u5_mult_82_CARRYB_5__12_, u5_mult_82_CARRYB_5__13_,
         u5_mult_82_CARRYB_5__14_, u5_mult_82_CARRYB_5__15_,
         u5_mult_82_CARRYB_5__16_, u5_mult_82_CARRYB_5__17_,
         u5_mult_82_CARRYB_5__18_, u5_mult_82_CARRYB_5__19_,
         u5_mult_82_CARRYB_5__20_, u5_mult_82_CARRYB_5__21_,
         u5_mult_82_CARRYB_5__22_, u5_mult_82_CARRYB_5__23_,
         u5_mult_82_CARRYB_5__24_, u5_mult_82_CARRYB_5__25_,
         u5_mult_82_CARRYB_5__26_, u5_mult_82_CARRYB_5__27_,
         u5_mult_82_CARRYB_5__28_, u5_mult_82_CARRYB_5__29_,
         u5_mult_82_CARRYB_5__30_, u5_mult_82_CARRYB_5__31_,
         u5_mult_82_CARRYB_5__32_, u5_mult_82_CARRYB_5__33_,
         u5_mult_82_CARRYB_5__34_, u5_mult_82_CARRYB_5__35_,
         u5_mult_82_CARRYB_5__36_, u5_mult_82_CARRYB_5__37_,
         u5_mult_82_CARRYB_5__38_, u5_mult_82_CARRYB_5__39_,
         u5_mult_82_CARRYB_5__40_, u5_mult_82_CARRYB_5__41_,
         u5_mult_82_CARRYB_5__42_, u5_mult_82_CARRYB_5__43_,
         u5_mult_82_CARRYB_5__44_, u5_mult_82_CARRYB_5__45_,
         u5_mult_82_CARRYB_5__46_, u5_mult_82_CARRYB_5__47_,
         u5_mult_82_CARRYB_5__48_, u5_mult_82_CARRYB_5__49_,
         u5_mult_82_CARRYB_5__50_, u5_mult_82_CARRYB_5__51_,
         u5_mult_82_CARRYB_6__0_, u5_mult_82_CARRYB_6__1_,
         u5_mult_82_CARRYB_6__2_, u5_mult_82_CARRYB_6__3_,
         u5_mult_82_CARRYB_6__4_, u5_mult_82_CARRYB_6__5_,
         u5_mult_82_CARRYB_6__6_, u5_mult_82_CARRYB_6__7_,
         u5_mult_82_CARRYB_6__8_, u5_mult_82_CARRYB_6__9_,
         u5_mult_82_CARRYB_6__10_, u5_mult_82_CARRYB_6__11_,
         u5_mult_82_CARRYB_6__12_, u5_mult_82_CARRYB_6__13_,
         u5_mult_82_CARRYB_6__14_, u5_mult_82_CARRYB_6__15_,
         u5_mult_82_CARRYB_6__16_, u5_mult_82_CARRYB_6__17_,
         u5_mult_82_CARRYB_6__18_, u5_mult_82_CARRYB_6__19_,
         u5_mult_82_CARRYB_6__20_, u5_mult_82_CARRYB_6__21_,
         u5_mult_82_CARRYB_6__22_, u5_mult_82_CARRYB_6__23_,
         u5_mult_82_CARRYB_6__24_, u5_mult_82_CARRYB_6__25_,
         u5_mult_82_CARRYB_6__26_, u5_mult_82_CARRYB_6__27_,
         u5_mult_82_CARRYB_6__28_, u5_mult_82_CARRYB_6__29_,
         u5_mult_82_CARRYB_6__30_, u5_mult_82_CARRYB_6__31_,
         u5_mult_82_CARRYB_6__32_, u5_mult_82_CARRYB_6__33_,
         u5_mult_82_CARRYB_6__34_, u5_mult_82_CARRYB_6__35_,
         u5_mult_82_CARRYB_6__36_, u5_mult_82_CARRYB_6__37_,
         u5_mult_82_CARRYB_6__38_, u5_mult_82_CARRYB_6__39_,
         u5_mult_82_CARRYB_6__40_, u5_mult_82_CARRYB_6__41_,
         u5_mult_82_CARRYB_6__42_, u5_mult_82_CARRYB_6__43_,
         u5_mult_82_CARRYB_6__44_, u5_mult_82_CARRYB_6__45_,
         u5_mult_82_CARRYB_6__46_, u5_mult_82_CARRYB_6__47_,
         u5_mult_82_CARRYB_6__48_, u5_mult_82_CARRYB_6__49_,
         u5_mult_82_CARRYB_6__50_, u5_mult_82_CARRYB_6__51_,
         u5_mult_82_CARRYB_7__0_, u5_mult_82_CARRYB_7__1_,
         u5_mult_82_CARRYB_7__2_, u5_mult_82_CARRYB_7__3_,
         u5_mult_82_CARRYB_7__4_, u5_mult_82_CARRYB_7__5_,
         u5_mult_82_CARRYB_7__6_, u5_mult_82_CARRYB_7__7_,
         u5_mult_82_CARRYB_7__8_, u5_mult_82_CARRYB_7__9_,
         u5_mult_82_CARRYB_7__10_, u5_mult_82_CARRYB_7__11_,
         u5_mult_82_CARRYB_7__12_, u5_mult_82_CARRYB_7__13_,
         u5_mult_82_CARRYB_7__14_, u5_mult_82_CARRYB_7__15_,
         u5_mult_82_CARRYB_7__16_, u5_mult_82_CARRYB_7__17_,
         u5_mult_82_CARRYB_7__18_, u5_mult_82_CARRYB_7__19_,
         u5_mult_82_CARRYB_7__20_, u5_mult_82_CARRYB_7__21_,
         u5_mult_82_CARRYB_7__22_, u5_mult_82_CARRYB_7__23_,
         u5_mult_82_CARRYB_7__24_, u5_mult_82_CARRYB_7__25_,
         u5_mult_82_CARRYB_7__26_, u5_mult_82_CARRYB_7__27_,
         u5_mult_82_CARRYB_7__28_, u5_mult_82_CARRYB_7__29_,
         u5_mult_82_CARRYB_7__30_, u5_mult_82_CARRYB_7__31_,
         u5_mult_82_CARRYB_7__32_, u5_mult_82_CARRYB_7__33_,
         u5_mult_82_CARRYB_7__34_, u5_mult_82_CARRYB_7__35_,
         u5_mult_82_CARRYB_7__36_, u5_mult_82_CARRYB_7__37_,
         u5_mult_82_CARRYB_7__38_, u5_mult_82_CARRYB_7__39_,
         u5_mult_82_CARRYB_7__40_, u5_mult_82_CARRYB_7__41_,
         u5_mult_82_CARRYB_7__42_, u5_mult_82_CARRYB_7__43_,
         u5_mult_82_CARRYB_7__44_, u5_mult_82_CARRYB_7__45_,
         u5_mult_82_CARRYB_7__46_, u5_mult_82_CARRYB_7__47_,
         u5_mult_82_CARRYB_7__48_, u5_mult_82_CARRYB_7__49_,
         u5_mult_82_CARRYB_7__50_, u5_mult_82_CARRYB_7__51_,
         u5_mult_82_CARRYB_8__0_, u5_mult_82_CARRYB_8__1_,
         u5_mult_82_CARRYB_8__2_, u5_mult_82_CARRYB_8__3_,
         u5_mult_82_CARRYB_8__4_, u5_mult_82_CARRYB_8__5_,
         u5_mult_82_CARRYB_8__6_, u5_mult_82_CARRYB_8__7_,
         u5_mult_82_CARRYB_8__8_, u5_mult_82_CARRYB_8__9_,
         u5_mult_82_CARRYB_8__10_, u5_mult_82_CARRYB_8__11_,
         u5_mult_82_CARRYB_8__12_, u5_mult_82_CARRYB_8__13_,
         u5_mult_82_CARRYB_8__14_, u5_mult_82_CARRYB_8__15_,
         u5_mult_82_CARRYB_8__16_, u5_mult_82_CARRYB_8__17_,
         u5_mult_82_CARRYB_8__18_, u5_mult_82_CARRYB_8__19_,
         u5_mult_82_CARRYB_8__20_, u5_mult_82_CARRYB_8__21_,
         u5_mult_82_CARRYB_8__22_, u5_mult_82_CARRYB_8__23_,
         u5_mult_82_CARRYB_8__24_, u5_mult_82_CARRYB_8__25_,
         u5_mult_82_CARRYB_8__26_, u5_mult_82_CARRYB_8__27_,
         u5_mult_82_CARRYB_8__28_, u5_mult_82_CARRYB_8__29_,
         u5_mult_82_CARRYB_8__30_, u5_mult_82_CARRYB_8__31_,
         u5_mult_82_CARRYB_8__32_, u5_mult_82_CARRYB_8__33_,
         u5_mult_82_CARRYB_8__34_, u5_mult_82_CARRYB_8__35_,
         u5_mult_82_CARRYB_8__36_, u5_mult_82_CARRYB_8__37_,
         u5_mult_82_CARRYB_8__38_, u5_mult_82_CARRYB_8__39_,
         u5_mult_82_CARRYB_8__40_, u5_mult_82_CARRYB_8__41_,
         u5_mult_82_CARRYB_8__42_, u5_mult_82_CARRYB_8__43_,
         u5_mult_82_CARRYB_8__44_, u5_mult_82_CARRYB_8__45_,
         u5_mult_82_CARRYB_8__46_, u5_mult_82_CARRYB_8__47_,
         u5_mult_82_CARRYB_8__48_, u5_mult_82_CARRYB_8__49_,
         u5_mult_82_CARRYB_8__50_, u5_mult_82_CARRYB_8__51_,
         u5_mult_82_CARRYB_9__0_, u5_mult_82_CARRYB_9__1_,
         u5_mult_82_CARRYB_9__2_, u5_mult_82_CARRYB_9__3_,
         u5_mult_82_CARRYB_9__4_, u5_mult_82_CARRYB_9__5_,
         u5_mult_82_CARRYB_9__6_, u5_mult_82_CARRYB_9__7_,
         u5_mult_82_CARRYB_9__8_, u5_mult_82_CARRYB_9__9_,
         u5_mult_82_CARRYB_9__10_, u5_mult_82_CARRYB_9__11_,
         u5_mult_82_CARRYB_9__12_, u5_mult_82_CARRYB_9__13_,
         u5_mult_82_CARRYB_9__14_, u5_mult_82_CARRYB_9__15_,
         u5_mult_82_CARRYB_9__16_, u5_mult_82_CARRYB_9__17_,
         u5_mult_82_CARRYB_9__18_, u5_mult_82_CARRYB_9__19_,
         u5_mult_82_CARRYB_9__20_, u5_mult_82_CARRYB_9__21_,
         u5_mult_82_CARRYB_9__22_, u5_mult_82_CARRYB_9__23_,
         u5_mult_82_CARRYB_9__24_, u5_mult_82_CARRYB_9__25_,
         u5_mult_82_CARRYB_9__26_, u5_mult_82_CARRYB_9__27_,
         u5_mult_82_CARRYB_9__28_, u5_mult_82_CARRYB_9__29_,
         u5_mult_82_CARRYB_9__30_, u5_mult_82_CARRYB_9__31_,
         u5_mult_82_CARRYB_9__32_, u5_mult_82_CARRYB_9__33_,
         u5_mult_82_CARRYB_9__34_, u5_mult_82_CARRYB_9__35_,
         u5_mult_82_CARRYB_9__36_, u5_mult_82_CARRYB_9__37_,
         u5_mult_82_CARRYB_9__38_, u5_mult_82_CARRYB_9__39_,
         u5_mult_82_CARRYB_9__40_, u5_mult_82_CARRYB_9__41_,
         u5_mult_82_CARRYB_9__42_, u5_mult_82_CARRYB_9__43_,
         u5_mult_82_CARRYB_9__44_, u5_mult_82_CARRYB_9__45_,
         u5_mult_82_CARRYB_9__46_, u5_mult_82_CARRYB_9__47_,
         u5_mult_82_CARRYB_9__48_, u5_mult_82_CARRYB_9__49_,
         u5_mult_82_CARRYB_9__50_, u5_mult_82_CARRYB_9__51_,
         u5_mult_82_CARRYB_10__0_, u5_mult_82_CARRYB_10__1_,
         u5_mult_82_CARRYB_10__2_, u5_mult_82_CARRYB_10__3_,
         u5_mult_82_CARRYB_10__4_, u5_mult_82_CARRYB_10__5_,
         u5_mult_82_CARRYB_10__6_, u5_mult_82_CARRYB_10__7_,
         u5_mult_82_CARRYB_10__8_, u5_mult_82_CARRYB_10__9_,
         u5_mult_82_CARRYB_10__10_, u5_mult_82_CARRYB_10__11_,
         u5_mult_82_CARRYB_10__12_, u5_mult_82_CARRYB_10__13_,
         u5_mult_82_CARRYB_10__14_, u5_mult_82_CARRYB_10__15_,
         u5_mult_82_CARRYB_10__16_, u5_mult_82_CARRYB_10__17_,
         u5_mult_82_CARRYB_10__18_, u5_mult_82_CARRYB_10__19_,
         u5_mult_82_CARRYB_10__20_, u5_mult_82_CARRYB_10__21_,
         u5_mult_82_CARRYB_10__22_, u5_mult_82_CARRYB_10__23_,
         u5_mult_82_CARRYB_10__24_, u5_mult_82_CARRYB_10__25_,
         u5_mult_82_CARRYB_10__26_, u5_mult_82_CARRYB_10__27_,
         u5_mult_82_CARRYB_10__28_, u5_mult_82_CARRYB_10__29_,
         u5_mult_82_CARRYB_10__30_, u5_mult_82_CARRYB_10__31_,
         u5_mult_82_CARRYB_10__32_, u5_mult_82_CARRYB_10__33_,
         u5_mult_82_CARRYB_10__34_, u5_mult_82_CARRYB_10__35_,
         u5_mult_82_CARRYB_10__36_, u5_mult_82_CARRYB_10__37_,
         u5_mult_82_CARRYB_10__38_, u5_mult_82_CARRYB_10__39_,
         u5_mult_82_CARRYB_10__40_, u5_mult_82_CARRYB_10__41_,
         u5_mult_82_CARRYB_10__42_, u5_mult_82_CARRYB_10__43_,
         u5_mult_82_CARRYB_10__44_, u5_mult_82_CARRYB_10__45_,
         u5_mult_82_CARRYB_10__46_, u5_mult_82_CARRYB_10__47_,
         u5_mult_82_CARRYB_10__48_, u5_mult_82_CARRYB_10__49_,
         u5_mult_82_CARRYB_10__50_, u5_mult_82_CARRYB_10__51_,
         u5_mult_82_CARRYB_11__0_, u5_mult_82_CARRYB_11__1_,
         u5_mult_82_CARRYB_11__2_, u5_mult_82_CARRYB_11__3_,
         u5_mult_82_CARRYB_11__4_, u5_mult_82_CARRYB_11__5_,
         u5_mult_82_CARRYB_11__6_, u5_mult_82_CARRYB_11__7_,
         u5_mult_82_CARRYB_11__8_, u5_mult_82_CARRYB_11__9_,
         u5_mult_82_CARRYB_11__10_, u5_mult_82_CARRYB_11__11_,
         u5_mult_82_CARRYB_11__12_, u5_mult_82_CARRYB_11__13_,
         u5_mult_82_CARRYB_11__14_, u5_mult_82_CARRYB_11__15_,
         u5_mult_82_CARRYB_11__16_, u5_mult_82_CARRYB_11__17_,
         u5_mult_82_CARRYB_11__18_, u5_mult_82_CARRYB_11__19_,
         u5_mult_82_CARRYB_11__20_, u5_mult_82_CARRYB_11__21_,
         u5_mult_82_CARRYB_11__22_, u5_mult_82_CARRYB_11__23_,
         u5_mult_82_CARRYB_11__24_, u5_mult_82_CARRYB_11__25_,
         u5_mult_82_CARRYB_11__26_, u5_mult_82_CARRYB_11__27_,
         u5_mult_82_CARRYB_11__28_, u5_mult_82_CARRYB_11__29_,
         u5_mult_82_CARRYB_11__30_, u5_mult_82_CARRYB_11__31_,
         u5_mult_82_CARRYB_11__32_, u5_mult_82_CARRYB_11__33_,
         u5_mult_82_CARRYB_11__34_, u5_mult_82_CARRYB_11__35_,
         u5_mult_82_CARRYB_11__36_, u5_mult_82_CARRYB_11__37_,
         u5_mult_82_CARRYB_11__38_, u5_mult_82_CARRYB_11__39_,
         u5_mult_82_CARRYB_11__40_, u5_mult_82_CARRYB_11__41_,
         u5_mult_82_CARRYB_11__42_, u5_mult_82_CARRYB_11__43_,
         u5_mult_82_CARRYB_11__44_, u5_mult_82_CARRYB_11__45_,
         u5_mult_82_CARRYB_11__46_, u5_mult_82_CARRYB_11__47_,
         u5_mult_82_CARRYB_11__48_, u5_mult_82_CARRYB_11__49_,
         u5_mult_82_CARRYB_11__50_, u5_mult_82_CARRYB_11__51_,
         u5_mult_82_CARRYB_12__0_, u5_mult_82_CARRYB_12__1_,
         u5_mult_82_CARRYB_12__2_, u5_mult_82_CARRYB_12__3_,
         u5_mult_82_CARRYB_12__4_, u5_mult_82_CARRYB_12__5_,
         u5_mult_82_CARRYB_12__6_, u5_mult_82_CARRYB_12__7_,
         u5_mult_82_CARRYB_12__8_, u5_mult_82_CARRYB_12__9_,
         u5_mult_82_CARRYB_12__10_, u5_mult_82_CARRYB_12__11_,
         u5_mult_82_CARRYB_12__12_, u5_mult_82_CARRYB_12__13_,
         u5_mult_82_CARRYB_12__14_, u5_mult_82_CARRYB_12__15_,
         u5_mult_82_CARRYB_12__16_, u5_mult_82_CARRYB_12__17_,
         u5_mult_82_CARRYB_12__18_, u5_mult_82_CARRYB_12__19_,
         u5_mult_82_CARRYB_12__20_, u5_mult_82_CARRYB_12__21_,
         u5_mult_82_CARRYB_12__22_, u5_mult_82_CARRYB_12__23_,
         u5_mult_82_CARRYB_12__24_, u5_mult_82_CARRYB_12__25_,
         u5_mult_82_CARRYB_12__26_, u5_mult_82_CARRYB_12__27_,
         u5_mult_82_CARRYB_12__28_, u5_mult_82_CARRYB_12__29_,
         u5_mult_82_CARRYB_12__30_, u5_mult_82_CARRYB_12__31_,
         u5_mult_82_CARRYB_12__32_, u5_mult_82_CARRYB_12__33_,
         u5_mult_82_CARRYB_12__34_, u5_mult_82_CARRYB_12__35_,
         u5_mult_82_CARRYB_12__36_, u5_mult_82_CARRYB_12__37_,
         u5_mult_82_CARRYB_12__38_, u5_mult_82_CARRYB_12__39_,
         u5_mult_82_CARRYB_12__40_, u5_mult_82_CARRYB_12__41_,
         u5_mult_82_CARRYB_12__42_, u5_mult_82_CARRYB_12__43_,
         u5_mult_82_CARRYB_12__44_, u5_mult_82_CARRYB_12__45_,
         u5_mult_82_CARRYB_12__46_, u5_mult_82_CARRYB_12__47_,
         u5_mult_82_CARRYB_12__48_, u5_mult_82_CARRYB_12__49_,
         u5_mult_82_CARRYB_12__50_, u5_mult_82_CARRYB_12__51_,
         u5_mult_82_CARRYB_13__0_, u5_mult_82_CARRYB_13__1_,
         u5_mult_82_CARRYB_13__2_, u5_mult_82_CARRYB_13__3_,
         u5_mult_82_CARRYB_13__4_, u5_mult_82_CARRYB_13__5_,
         u5_mult_82_CARRYB_13__6_, u5_mult_82_CARRYB_13__7_,
         u5_mult_82_CARRYB_13__8_, u5_mult_82_CARRYB_13__9_,
         u5_mult_82_CARRYB_13__10_, u5_mult_82_CARRYB_13__11_,
         u5_mult_82_CARRYB_13__12_, u5_mult_82_CARRYB_13__13_,
         u5_mult_82_CARRYB_13__14_, u5_mult_82_CARRYB_13__15_,
         u5_mult_82_CARRYB_13__16_, u5_mult_82_CARRYB_13__17_,
         u5_mult_82_CARRYB_13__18_, u5_mult_82_CARRYB_13__19_,
         u5_mult_82_CARRYB_13__20_, u5_mult_82_CARRYB_13__21_,
         u5_mult_82_CARRYB_13__22_, u5_mult_82_CARRYB_13__23_,
         u5_mult_82_CARRYB_13__24_, u5_mult_82_CARRYB_13__25_,
         u5_mult_82_CARRYB_13__26_, u5_mult_82_CARRYB_13__27_,
         u5_mult_82_CARRYB_13__28_, u5_mult_82_CARRYB_13__29_,
         u5_mult_82_CARRYB_13__30_, u5_mult_82_CARRYB_13__31_,
         u5_mult_82_CARRYB_13__32_, u5_mult_82_CARRYB_13__33_,
         u5_mult_82_CARRYB_13__34_, u5_mult_82_CARRYB_13__35_,
         u5_mult_82_CARRYB_13__36_, u5_mult_82_CARRYB_13__37_,
         u5_mult_82_CARRYB_13__38_, u5_mult_82_CARRYB_13__39_,
         u5_mult_82_CARRYB_13__40_, u5_mult_82_CARRYB_13__41_,
         u5_mult_82_CARRYB_13__42_, u5_mult_82_CARRYB_13__43_,
         u5_mult_82_CARRYB_13__44_, u5_mult_82_CARRYB_13__45_,
         u5_mult_82_CARRYB_13__46_, u5_mult_82_CARRYB_13__47_,
         u5_mult_82_CARRYB_13__48_, u5_mult_82_CARRYB_13__49_,
         u5_mult_82_CARRYB_13__50_, u5_mult_82_CARRYB_13__51_,
         u5_mult_82_CARRYB_14__0_, u5_mult_82_CARRYB_14__1_,
         u5_mult_82_CARRYB_14__2_, u5_mult_82_CARRYB_14__3_,
         u5_mult_82_CARRYB_14__4_, u5_mult_82_CARRYB_14__5_,
         u5_mult_82_CARRYB_14__6_, u5_mult_82_CARRYB_14__7_,
         u5_mult_82_CARRYB_14__8_, u5_mult_82_CARRYB_14__9_,
         u5_mult_82_CARRYB_14__10_, u5_mult_82_CARRYB_14__11_,
         u5_mult_82_CARRYB_14__12_, u5_mult_82_CARRYB_14__13_,
         u5_mult_82_CARRYB_14__14_, u5_mult_82_CARRYB_14__15_,
         u5_mult_82_CARRYB_14__16_, u5_mult_82_CARRYB_14__17_,
         u5_mult_82_CARRYB_14__18_, u5_mult_82_SUMB_2__1_,
         u5_mult_82_SUMB_2__2_, u5_mult_82_SUMB_2__3_, u5_mult_82_SUMB_2__4_,
         u5_mult_82_SUMB_2__5_, u5_mult_82_SUMB_2__6_, u5_mult_82_SUMB_2__7_,
         u5_mult_82_SUMB_2__8_, u5_mult_82_SUMB_2__9_, u5_mult_82_SUMB_2__10_,
         u5_mult_82_SUMB_2__11_, u5_mult_82_SUMB_2__12_,
         u5_mult_82_SUMB_2__13_, u5_mult_82_SUMB_2__14_,
         u5_mult_82_SUMB_2__15_, u5_mult_82_SUMB_2__16_,
         u5_mult_82_SUMB_2__17_, u5_mult_82_SUMB_2__18_,
         u5_mult_82_SUMB_2__19_, u5_mult_82_SUMB_2__20_,
         u5_mult_82_SUMB_2__21_, u5_mult_82_SUMB_2__22_,
         u5_mult_82_SUMB_2__23_, u5_mult_82_SUMB_2__24_,
         u5_mult_82_SUMB_2__25_, u5_mult_82_SUMB_2__26_,
         u5_mult_82_SUMB_2__27_, u5_mult_82_SUMB_2__28_,
         u5_mult_82_SUMB_2__29_, u5_mult_82_SUMB_2__30_,
         u5_mult_82_SUMB_2__31_, u5_mult_82_SUMB_2__32_,
         u5_mult_82_SUMB_2__33_, u5_mult_82_SUMB_2__34_,
         u5_mult_82_SUMB_2__35_, u5_mult_82_SUMB_2__36_,
         u5_mult_82_SUMB_2__37_, u5_mult_82_SUMB_2__38_,
         u5_mult_82_SUMB_2__39_, u5_mult_82_SUMB_2__40_,
         u5_mult_82_SUMB_2__41_, u5_mult_82_SUMB_2__42_,
         u5_mult_82_SUMB_2__43_, u5_mult_82_SUMB_2__44_,
         u5_mult_82_SUMB_2__45_, u5_mult_82_SUMB_2__46_,
         u5_mult_82_SUMB_2__47_, u5_mult_82_SUMB_2__48_,
         u5_mult_82_SUMB_2__49_, u5_mult_82_SUMB_2__50_,
         u5_mult_82_SUMB_2__51_, u5_mult_82_SUMB_3__1_, u5_mult_82_SUMB_3__2_,
         u5_mult_82_SUMB_3__3_, u5_mult_82_SUMB_3__4_, u5_mult_82_SUMB_3__5_,
         u5_mult_82_SUMB_3__6_, u5_mult_82_SUMB_3__7_, u5_mult_82_SUMB_3__8_,
         u5_mult_82_SUMB_3__9_, u5_mult_82_SUMB_3__10_, u5_mult_82_SUMB_3__11_,
         u5_mult_82_SUMB_3__12_, u5_mult_82_SUMB_3__13_,
         u5_mult_82_SUMB_3__14_, u5_mult_82_SUMB_3__15_,
         u5_mult_82_SUMB_3__16_, u5_mult_82_SUMB_3__17_,
         u5_mult_82_SUMB_3__18_, u5_mult_82_SUMB_3__19_,
         u5_mult_82_SUMB_3__20_, u5_mult_82_SUMB_3__21_,
         u5_mult_82_SUMB_3__22_, u5_mult_82_SUMB_3__23_,
         u5_mult_82_SUMB_3__24_, u5_mult_82_SUMB_3__25_,
         u5_mult_82_SUMB_3__26_, u5_mult_82_SUMB_3__27_,
         u5_mult_82_SUMB_3__28_, u5_mult_82_SUMB_3__29_,
         u5_mult_82_SUMB_3__30_, u5_mult_82_SUMB_3__31_,
         u5_mult_82_SUMB_3__32_, u5_mult_82_SUMB_3__33_,
         u5_mult_82_SUMB_3__34_, u5_mult_82_SUMB_3__35_,
         u5_mult_82_SUMB_3__36_, u5_mult_82_SUMB_3__37_,
         u5_mult_82_SUMB_3__38_, u5_mult_82_SUMB_3__39_,
         u5_mult_82_SUMB_3__40_, u5_mult_82_SUMB_3__41_,
         u5_mult_82_SUMB_3__42_, u5_mult_82_SUMB_3__43_,
         u5_mult_82_SUMB_3__44_, u5_mult_82_SUMB_3__45_,
         u5_mult_82_SUMB_3__46_, u5_mult_82_SUMB_3__47_,
         u5_mult_82_SUMB_3__48_, u5_mult_82_SUMB_3__49_,
         u5_mult_82_SUMB_3__50_, u5_mult_82_SUMB_3__51_, u5_mult_82_SUMB_4__1_,
         u5_mult_82_SUMB_4__2_, u5_mult_82_SUMB_4__3_, u5_mult_82_SUMB_4__4_,
         u5_mult_82_SUMB_4__5_, u5_mult_82_SUMB_4__6_, u5_mult_82_SUMB_4__7_,
         u5_mult_82_SUMB_4__8_, u5_mult_82_SUMB_4__9_, u5_mult_82_SUMB_4__10_,
         u5_mult_82_SUMB_4__11_, u5_mult_82_SUMB_4__12_,
         u5_mult_82_SUMB_4__13_, u5_mult_82_SUMB_4__14_,
         u5_mult_82_SUMB_4__15_, u5_mult_82_SUMB_4__16_,
         u5_mult_82_SUMB_4__17_, u5_mult_82_SUMB_4__18_,
         u5_mult_82_SUMB_4__19_, u5_mult_82_SUMB_4__20_,
         u5_mult_82_SUMB_4__21_, u5_mult_82_SUMB_4__22_,
         u5_mult_82_SUMB_4__23_, u5_mult_82_SUMB_4__24_,
         u5_mult_82_SUMB_4__25_, u5_mult_82_SUMB_4__26_,
         u5_mult_82_SUMB_4__27_, u5_mult_82_SUMB_4__28_,
         u5_mult_82_SUMB_4__29_, u5_mult_82_SUMB_4__30_,
         u5_mult_82_SUMB_4__31_, u5_mult_82_SUMB_4__32_,
         u5_mult_82_SUMB_4__33_, u5_mult_82_SUMB_4__34_,
         u5_mult_82_SUMB_4__35_, u5_mult_82_SUMB_4__36_,
         u5_mult_82_CARRYB_2__0_, u5_mult_82_CARRYB_2__1_,
         u5_mult_82_CARRYB_2__2_, u5_mult_82_CARRYB_2__3_,
         u5_mult_82_CARRYB_2__4_, u5_mult_82_CARRYB_2__5_,
         u5_mult_82_CARRYB_2__6_, u5_mult_82_CARRYB_2__7_,
         u5_mult_82_CARRYB_2__8_, u5_mult_82_CARRYB_2__9_,
         u5_mult_82_CARRYB_2__10_, u5_mult_82_CARRYB_2__11_,
         u5_mult_82_CARRYB_2__12_, u5_mult_82_CARRYB_2__13_,
         u5_mult_82_CARRYB_2__14_, u5_mult_82_CARRYB_2__15_,
         u5_mult_82_CARRYB_2__16_, u5_mult_82_CARRYB_2__17_,
         u5_mult_82_CARRYB_2__18_, u5_mult_82_CARRYB_2__19_,
         u5_mult_82_CARRYB_2__20_, u5_mult_82_CARRYB_2__21_,
         u5_mult_82_CARRYB_2__22_, u5_mult_82_CARRYB_2__23_,
         u5_mult_82_CARRYB_2__24_, u5_mult_82_CARRYB_2__25_,
         u5_mult_82_CARRYB_2__26_, u5_mult_82_CARRYB_2__27_,
         u5_mult_82_CARRYB_2__28_, u5_mult_82_CARRYB_2__29_,
         u5_mult_82_CARRYB_2__30_, u5_mult_82_CARRYB_2__31_,
         u5_mult_82_CARRYB_2__32_, u5_mult_82_CARRYB_2__33_,
         u5_mult_82_CARRYB_2__34_, u5_mult_82_CARRYB_2__35_,
         u5_mult_82_CARRYB_2__36_, u5_mult_82_CARRYB_2__37_,
         u5_mult_82_CARRYB_2__38_, u5_mult_82_CARRYB_2__39_,
         u5_mult_82_CARRYB_2__40_, u5_mult_82_CARRYB_2__41_,
         u5_mult_82_CARRYB_2__42_, u5_mult_82_CARRYB_2__43_,
         u5_mult_82_CARRYB_2__44_, u5_mult_82_CARRYB_2__45_,
         u5_mult_82_CARRYB_2__46_, u5_mult_82_CARRYB_2__47_,
         u5_mult_82_CARRYB_2__48_, u5_mult_82_CARRYB_2__49_,
         u5_mult_82_CARRYB_2__50_, u5_mult_82_CARRYB_2__51_,
         u5_mult_82_CARRYB_3__0_, u5_mult_82_CARRYB_3__1_,
         u5_mult_82_CARRYB_3__2_, u5_mult_82_CARRYB_3__3_,
         u5_mult_82_CARRYB_3__4_, u5_mult_82_CARRYB_3__5_,
         u5_mult_82_CARRYB_3__6_, u5_mult_82_CARRYB_3__7_,
         u5_mult_82_CARRYB_3__8_, u5_mult_82_CARRYB_3__9_,
         u5_mult_82_CARRYB_3__10_, u5_mult_82_CARRYB_3__11_,
         u5_mult_82_CARRYB_3__12_, u5_mult_82_CARRYB_3__13_,
         u5_mult_82_CARRYB_3__14_, u5_mult_82_CARRYB_3__15_,
         u5_mult_82_CARRYB_3__16_, u5_mult_82_CARRYB_3__17_,
         u5_mult_82_CARRYB_3__18_, u5_mult_82_CARRYB_3__19_,
         u5_mult_82_CARRYB_3__20_, u5_mult_82_CARRYB_3__21_,
         u5_mult_82_CARRYB_3__22_, u5_mult_82_CARRYB_3__23_,
         u5_mult_82_CARRYB_3__24_, u5_mult_82_CARRYB_3__25_,
         u5_mult_82_CARRYB_3__26_, u5_mult_82_CARRYB_3__27_,
         u5_mult_82_CARRYB_3__28_, u5_mult_82_CARRYB_3__29_,
         u5_mult_82_CARRYB_3__30_, u5_mult_82_CARRYB_3__31_,
         u5_mult_82_CARRYB_3__32_, u5_mult_82_CARRYB_3__33_,
         u5_mult_82_CARRYB_3__34_, u5_mult_82_CARRYB_3__35_,
         u5_mult_82_CARRYB_3__36_, u5_mult_82_CARRYB_3__37_,
         u5_mult_82_CARRYB_3__38_, u5_mult_82_CARRYB_3__39_,
         u5_mult_82_CARRYB_3__40_, u5_mult_82_CARRYB_3__41_,
         u5_mult_82_CARRYB_3__42_, u5_mult_82_CARRYB_3__43_,
         u5_mult_82_CARRYB_3__44_, u5_mult_82_CARRYB_3__45_,
         u5_mult_82_CARRYB_3__46_, u5_mult_82_CARRYB_3__47_,
         u5_mult_82_CARRYB_3__48_, u5_mult_82_CARRYB_3__49_,
         u5_mult_82_CARRYB_3__50_, u5_mult_82_CARRYB_3__51_,
         u5_mult_82_CARRYB_4__0_, u5_mult_82_CARRYB_4__1_,
         u5_mult_82_CARRYB_4__2_, u5_mult_82_CARRYB_4__3_,
         u5_mult_82_CARRYB_4__4_, u5_mult_82_CARRYB_4__5_,
         u5_mult_82_CARRYB_4__6_, u5_mult_82_CARRYB_4__7_,
         u5_mult_82_CARRYB_4__8_, u5_mult_82_CARRYB_4__9_,
         u5_mult_82_CARRYB_4__10_, u5_mult_82_CARRYB_4__11_,
         u5_mult_82_CARRYB_4__12_, u5_mult_82_CARRYB_4__13_,
         u5_mult_82_CARRYB_4__14_, u5_mult_82_CARRYB_4__15_,
         u5_mult_82_CARRYB_4__16_, u5_mult_82_CARRYB_4__17_,
         u5_mult_82_CARRYB_4__18_, u5_mult_82_CARRYB_4__19_,
         u5_mult_82_CARRYB_4__20_, u5_mult_82_CARRYB_4__21_,
         u5_mult_82_CARRYB_4__22_, u5_mult_82_CARRYB_4__23_,
         u5_mult_82_CARRYB_4__24_, u5_mult_82_CARRYB_4__25_,
         u5_mult_82_CARRYB_4__26_, u5_mult_82_CARRYB_4__27_,
         u5_mult_82_CARRYB_4__28_, u5_mult_82_CARRYB_4__29_,
         u5_mult_82_CARRYB_4__30_, u5_mult_82_CARRYB_4__31_,
         u5_mult_82_CARRYB_4__32_, u5_mult_82_CARRYB_4__33_,
         u5_mult_82_CARRYB_4__34_, u5_mult_82_CARRYB_4__35_,
         u5_mult_82_CARRYB_4__36_, u5_mult_82_ab_0__1_, u5_mult_82_ab_0__2_,
         u5_mult_82_ab_0__3_, u5_mult_82_ab_0__4_, u5_mult_82_ab_0__5_,
         u5_mult_82_ab_0__6_, u5_mult_82_ab_0__7_, u5_mult_82_ab_0__8_,
         u5_mult_82_ab_0__9_, u5_mult_82_ab_0__10_, u5_mult_82_ab_0__11_,
         u5_mult_82_ab_0__12_, u5_mult_82_ab_0__13_, u5_mult_82_ab_0__14_,
         u5_mult_82_ab_0__15_, u5_mult_82_ab_0__16_, u5_mult_82_ab_0__17_,
         u5_mult_82_ab_0__18_, u5_mult_82_ab_0__19_, u5_mult_82_ab_0__20_,
         u5_mult_82_ab_0__21_, u5_mult_82_ab_0__22_, u5_mult_82_ab_0__23_,
         u5_mult_82_ab_0__24_, u5_mult_82_ab_0__25_, u5_mult_82_ab_0__26_,
         u5_mult_82_ab_0__27_, u5_mult_82_ab_0__28_, u5_mult_82_ab_0__29_,
         u5_mult_82_ab_0__30_, u5_mult_82_ab_0__31_, u5_mult_82_ab_0__32_,
         u5_mult_82_ab_0__33_, u5_mult_82_ab_0__34_, u5_mult_82_ab_0__35_,
         u5_mult_82_ab_0__36_, u5_mult_82_ab_0__37_, u5_mult_82_ab_0__38_,
         u5_mult_82_ab_0__39_, u5_mult_82_ab_0__40_, u5_mult_82_ab_0__41_,
         u5_mult_82_ab_0__42_, u5_mult_82_ab_0__43_, u5_mult_82_ab_0__44_,
         u5_mult_82_ab_0__45_, u5_mult_82_ab_0__46_, u5_mult_82_ab_0__47_,
         u5_mult_82_ab_0__48_, u5_mult_82_ab_0__49_, u5_mult_82_ab_0__50_,
         u5_mult_82_ab_0__51_, u5_mult_82_ab_0__52_, u5_mult_82_ab_1__0_,
         u5_mult_82_ab_1__1_, u5_mult_82_ab_1__2_, u5_mult_82_ab_1__3_,
         u5_mult_82_ab_1__4_, u5_mult_82_ab_1__5_, u5_mult_82_ab_1__6_,
         u5_mult_82_ab_1__7_, u5_mult_82_ab_1__8_, u5_mult_82_ab_1__9_,
         u5_mult_82_ab_1__10_, u5_mult_82_ab_1__11_, u5_mult_82_ab_1__12_,
         u5_mult_82_ab_1__13_, u5_mult_82_ab_1__14_, u5_mult_82_ab_1__15_,
         u5_mult_82_ab_1__16_, u5_mult_82_ab_1__17_, u5_mult_82_ab_1__18_,
         u5_mult_82_ab_1__19_, u5_mult_82_ab_1__20_, u5_mult_82_ab_1__21_,
         u5_mult_82_ab_1__22_, u5_mult_82_ab_1__23_, u5_mult_82_ab_1__24_,
         u5_mult_82_ab_1__25_, u5_mult_82_ab_1__26_, u5_mult_82_ab_1__27_,
         u5_mult_82_ab_1__28_, u5_mult_82_ab_1__29_, u5_mult_82_ab_1__30_,
         u5_mult_82_ab_1__31_, u5_mult_82_ab_1__32_, u5_mult_82_ab_1__33_,
         u5_mult_82_ab_1__34_, u5_mult_82_ab_1__35_, u5_mult_82_ab_1__36_,
         u5_mult_82_ab_1__37_, u5_mult_82_ab_1__38_, u5_mult_82_ab_1__39_,
         u5_mult_82_ab_1__40_, u5_mult_82_ab_1__41_, u5_mult_82_ab_1__42_,
         u5_mult_82_ab_1__43_, u5_mult_82_ab_1__44_, u5_mult_82_ab_1__45_,
         u5_mult_82_ab_1__46_, u5_mult_82_ab_1__47_, u5_mult_82_ab_1__48_,
         u5_mult_82_ab_1__49_, u5_mult_82_ab_1__50_, u5_mult_82_ab_1__51_,
         u5_mult_82_ab_1__52_, u5_mult_82_ab_2__0_, u5_mult_82_ab_2__1_,
         u5_mult_82_ab_2__2_, u5_mult_82_ab_2__3_, u5_mult_82_ab_2__4_,
         u5_mult_82_ab_2__5_, u5_mult_82_ab_2__6_, u5_mult_82_ab_2__7_,
         u5_mult_82_ab_2__8_, u5_mult_82_ab_2__9_, u5_mult_82_ab_2__10_,
         u5_mult_82_ab_2__11_, u5_mult_82_ab_2__12_, u5_mult_82_ab_2__13_,
         u5_mult_82_ab_2__14_, u5_mult_82_ab_2__15_, u5_mult_82_ab_2__16_,
         u5_mult_82_ab_2__17_, u5_mult_82_ab_2__18_, u5_mult_82_ab_2__19_,
         u5_mult_82_ab_2__20_, u5_mult_82_ab_2__21_, u5_mult_82_ab_2__22_,
         u5_mult_82_ab_2__23_, u5_mult_82_ab_2__24_, u5_mult_82_ab_2__25_,
         u5_mult_82_ab_2__26_, u5_mult_82_ab_2__27_, u5_mult_82_ab_2__28_,
         u5_mult_82_ab_2__29_, u5_mult_82_ab_2__30_, u5_mult_82_ab_2__31_,
         u5_mult_82_ab_2__32_, u5_mult_82_ab_2__33_, u5_mult_82_ab_2__34_,
         u5_mult_82_ab_2__35_, u5_mult_82_ab_2__36_, u5_mult_82_ab_2__37_,
         u5_mult_82_ab_2__38_, u5_mult_82_ab_2__39_, u5_mult_82_ab_2__40_,
         u5_mult_82_ab_2__41_, u5_mult_82_ab_2__42_, u5_mult_82_ab_2__43_,
         u5_mult_82_ab_2__44_, u5_mult_82_ab_2__45_, u5_mult_82_ab_2__46_,
         u5_mult_82_ab_2__47_, u5_mult_82_ab_2__48_, u5_mult_82_ab_2__49_,
         u5_mult_82_ab_2__50_, u5_mult_82_ab_2__51_, u5_mult_82_ab_2__52_,
         u5_mult_82_ab_3__0_, u5_mult_82_ab_3__1_, u5_mult_82_ab_3__2_,
         u5_mult_82_ab_3__3_, u5_mult_82_ab_3__4_, u5_mult_82_ab_3__5_,
         u5_mult_82_ab_3__6_, u5_mult_82_ab_3__7_, u5_mult_82_ab_3__8_,
         u5_mult_82_ab_3__9_, u5_mult_82_ab_3__10_, u5_mult_82_ab_3__11_,
         u5_mult_82_ab_3__12_, u5_mult_82_ab_3__13_, u5_mult_82_ab_3__14_,
         u5_mult_82_ab_3__15_, u5_mult_82_ab_3__16_, u5_mult_82_ab_3__17_,
         u5_mult_82_ab_3__18_, u5_mult_82_ab_3__19_, u5_mult_82_ab_3__20_,
         u5_mult_82_ab_3__21_, u5_mult_82_ab_3__22_, u5_mult_82_ab_3__23_,
         u5_mult_82_ab_3__24_, u5_mult_82_ab_3__25_, u5_mult_82_ab_3__26_,
         u5_mult_82_ab_3__27_, u5_mult_82_ab_3__28_, u5_mult_82_ab_3__29_,
         u5_mult_82_ab_3__30_, u5_mult_82_ab_3__31_, u5_mult_82_ab_3__32_,
         u5_mult_82_ab_3__33_, u5_mult_82_ab_3__34_, u5_mult_82_ab_3__35_,
         u5_mult_82_ab_3__36_, u5_mult_82_ab_3__37_, u5_mult_82_ab_3__38_,
         u5_mult_82_ab_3__39_, u5_mult_82_ab_3__40_, u5_mult_82_ab_3__41_,
         u5_mult_82_ab_3__42_, u5_mult_82_ab_3__43_, u5_mult_82_ab_3__44_,
         u5_mult_82_ab_3__45_, u5_mult_82_ab_3__46_, u5_mult_82_ab_3__47_,
         u5_mult_82_ab_3__48_, u5_mult_82_ab_3__49_, u5_mult_82_ab_3__50_,
         u5_mult_82_ab_3__51_, u5_mult_82_ab_3__52_, u5_mult_82_ab_4__0_,
         u5_mult_82_ab_4__1_, u5_mult_82_ab_4__2_, u5_mult_82_ab_4__3_,
         u5_mult_82_ab_4__4_, u5_mult_82_ab_4__5_, u5_mult_82_ab_4__6_,
         u5_mult_82_ab_4__7_, u5_mult_82_ab_4__8_, u5_mult_82_ab_4__9_,
         u5_mult_82_ab_4__10_, u5_mult_82_ab_4__11_, u5_mult_82_ab_4__12_,
         u5_mult_82_ab_4__13_, u5_mult_82_ab_4__14_, u5_mult_82_ab_4__15_,
         u5_mult_82_ab_4__16_, u5_mult_82_ab_4__17_, u5_mult_82_ab_4__18_,
         u5_mult_82_ab_4__19_, u5_mult_82_ab_4__20_, u5_mult_82_ab_4__21_,
         u5_mult_82_ab_4__22_, u5_mult_82_ab_4__23_, u5_mult_82_ab_4__24_,
         u5_mult_82_ab_4__25_, u5_mult_82_ab_4__26_, u5_mult_82_ab_4__27_,
         u5_mult_82_ab_4__28_, u5_mult_82_ab_4__29_, u5_mult_82_ab_4__30_,
         u5_mult_82_ab_4__31_, u5_mult_82_ab_4__32_, u5_mult_82_ab_4__33_,
         u5_mult_82_ab_4__34_, u5_mult_82_ab_4__35_, u5_mult_82_ab_4__36_,
         u5_mult_82_ab_4__37_, u5_mult_82_ab_4__38_, u5_mult_82_ab_4__39_,
         u5_mult_82_ab_4__40_, u5_mult_82_ab_4__41_, u5_mult_82_ab_4__42_,
         u5_mult_82_ab_4__43_, u5_mult_82_ab_4__44_, u5_mult_82_ab_4__45_,
         u5_mult_82_ab_4__46_, u5_mult_82_ab_4__47_, u5_mult_82_ab_4__48_,
         u5_mult_82_ab_4__49_, u5_mult_82_ab_4__50_, u5_mult_82_ab_4__51_,
         u5_mult_82_ab_4__52_, u5_mult_82_ab_5__0_, u5_mult_82_ab_5__1_,
         u5_mult_82_ab_5__2_, u5_mult_82_ab_5__3_, u5_mult_82_ab_5__4_,
         u5_mult_82_ab_5__5_, u5_mult_82_ab_5__6_, u5_mult_82_ab_5__7_,
         u5_mult_82_ab_5__8_, u5_mult_82_ab_5__9_, u5_mult_82_ab_5__10_,
         u5_mult_82_ab_5__11_, u5_mult_82_ab_5__12_, u5_mult_82_ab_5__13_,
         u5_mult_82_ab_5__14_, u5_mult_82_ab_5__15_, u5_mult_82_ab_5__16_,
         u5_mult_82_ab_5__17_, u5_mult_82_ab_5__18_, u5_mult_82_ab_5__19_,
         u5_mult_82_ab_5__20_, u5_mult_82_ab_5__21_, u5_mult_82_ab_5__22_,
         u5_mult_82_ab_5__23_, u5_mult_82_ab_5__24_, u5_mult_82_ab_5__25_,
         u5_mult_82_ab_5__26_, u5_mult_82_ab_5__27_, u5_mult_82_ab_5__28_,
         u5_mult_82_ab_5__29_, u5_mult_82_ab_5__30_, u5_mult_82_ab_5__31_,
         u5_mult_82_ab_5__32_, u5_mult_82_ab_5__33_, u5_mult_82_ab_5__34_,
         u5_mult_82_ab_5__35_, u5_mult_82_ab_5__36_, u5_mult_82_ab_5__37_,
         u5_mult_82_ab_5__38_, u5_mult_82_ab_5__39_, u5_mult_82_ab_5__40_,
         u5_mult_82_ab_5__41_, u5_mult_82_ab_5__42_, u5_mult_82_ab_5__43_,
         u5_mult_82_ab_5__44_, u5_mult_82_ab_5__45_, u5_mult_82_ab_5__46_,
         u5_mult_82_ab_5__47_, u5_mult_82_ab_5__48_, u5_mult_82_ab_5__49_,
         u5_mult_82_ab_5__50_, u5_mult_82_ab_5__51_, u5_mult_82_ab_5__52_,
         u5_mult_82_ab_6__0_, u5_mult_82_ab_6__1_, u5_mult_82_ab_6__2_,
         u5_mult_82_ab_6__3_, u5_mult_82_ab_6__4_, u5_mult_82_ab_6__5_,
         u5_mult_82_ab_6__6_, u5_mult_82_ab_6__7_, u5_mult_82_ab_6__8_,
         u5_mult_82_ab_6__9_, u5_mult_82_ab_6__10_, u5_mult_82_ab_6__11_,
         u5_mult_82_ab_6__12_, u5_mult_82_ab_6__13_, u5_mult_82_ab_6__14_,
         u5_mult_82_ab_6__15_, u5_mult_82_ab_6__16_, u5_mult_82_ab_6__17_,
         u5_mult_82_ab_6__18_, u5_mult_82_ab_6__19_, u5_mult_82_ab_6__20_,
         u5_mult_82_ab_6__21_, u5_mult_82_ab_6__22_, u5_mult_82_ab_6__23_,
         u5_mult_82_ab_6__24_, u5_mult_82_ab_6__25_, u5_mult_82_ab_6__26_,
         u5_mult_82_ab_6__27_, u5_mult_82_ab_6__28_, u5_mult_82_ab_6__29_,
         u5_mult_82_ab_6__30_, u5_mult_82_ab_6__31_, u5_mult_82_ab_6__32_,
         u5_mult_82_ab_6__33_, u5_mult_82_ab_6__34_, u5_mult_82_ab_6__35_,
         u5_mult_82_ab_6__36_, u5_mult_82_ab_6__37_, u5_mult_82_ab_6__38_,
         u5_mult_82_ab_6__39_, u5_mult_82_ab_6__40_, u5_mult_82_ab_6__41_,
         u5_mult_82_ab_6__42_, u5_mult_82_ab_6__43_, u5_mult_82_ab_6__44_,
         u5_mult_82_ab_6__45_, u5_mult_82_ab_6__46_, u5_mult_82_ab_6__47_,
         u5_mult_82_ab_6__48_, u5_mult_82_ab_6__49_, u5_mult_82_ab_6__50_,
         u5_mult_82_ab_6__51_, u5_mult_82_ab_6__52_, u5_mult_82_ab_7__0_,
         u5_mult_82_ab_7__1_, u5_mult_82_ab_7__2_, u5_mult_82_ab_7__3_,
         u5_mult_82_ab_7__4_, u5_mult_82_ab_7__5_, u5_mult_82_ab_7__6_,
         u5_mult_82_ab_7__7_, u5_mult_82_ab_7__8_, u5_mult_82_ab_7__9_,
         u5_mult_82_ab_7__10_, u5_mult_82_ab_7__11_, u5_mult_82_ab_7__12_,
         u5_mult_82_ab_7__13_, u5_mult_82_ab_7__14_, u5_mult_82_ab_7__15_,
         u5_mult_82_ab_7__16_, u5_mult_82_ab_7__17_, u5_mult_82_ab_7__18_,
         u5_mult_82_ab_7__19_, u5_mult_82_ab_7__20_, u5_mult_82_ab_7__21_,
         u5_mult_82_ab_7__22_, u5_mult_82_ab_7__23_, u5_mult_82_ab_7__24_,
         u5_mult_82_ab_7__25_, u5_mult_82_ab_7__26_, u5_mult_82_ab_7__27_,
         u5_mult_82_ab_7__28_, u5_mult_82_ab_7__29_, u5_mult_82_ab_7__30_,
         u5_mult_82_ab_7__31_, u5_mult_82_ab_7__32_, u5_mult_82_ab_7__33_,
         u5_mult_82_ab_7__34_, u5_mult_82_ab_7__35_, u5_mult_82_ab_7__36_,
         u5_mult_82_ab_7__37_, u5_mult_82_ab_7__38_, u5_mult_82_ab_7__39_,
         u5_mult_82_ab_7__40_, u5_mult_82_ab_7__41_, u5_mult_82_ab_7__42_,
         u5_mult_82_ab_7__43_, u5_mult_82_ab_7__44_, u5_mult_82_ab_7__45_,
         u5_mult_82_ab_7__46_, u5_mult_82_ab_7__47_, u5_mult_82_ab_7__48_,
         u5_mult_82_ab_7__49_, u5_mult_82_ab_7__50_, u5_mult_82_ab_7__51_,
         u5_mult_82_ab_7__52_, u5_mult_82_ab_8__0_, u5_mult_82_ab_8__1_,
         u5_mult_82_ab_8__2_, u5_mult_82_ab_8__3_, u5_mult_82_ab_8__4_,
         u5_mult_82_ab_8__5_, u5_mult_82_ab_8__6_, u5_mult_82_ab_8__7_,
         u5_mult_82_ab_8__8_, u5_mult_82_ab_8__9_, u5_mult_82_ab_8__10_,
         u5_mult_82_ab_8__11_, u5_mult_82_ab_8__12_, u5_mult_82_ab_8__13_,
         u5_mult_82_ab_8__14_, u5_mult_82_ab_8__15_, u5_mult_82_ab_8__16_,
         u5_mult_82_ab_8__17_, u5_mult_82_ab_8__18_, u5_mult_82_ab_8__19_,
         u5_mult_82_ab_8__20_, u5_mult_82_ab_8__21_, u5_mult_82_ab_8__22_,
         u5_mult_82_ab_8__23_, u5_mult_82_ab_8__24_, u5_mult_82_ab_8__25_,
         u5_mult_82_ab_8__26_, u5_mult_82_ab_8__27_, u5_mult_82_ab_8__28_,
         u5_mult_82_ab_8__29_, u5_mult_82_ab_8__30_, u5_mult_82_ab_8__31_,
         u5_mult_82_ab_8__32_, u5_mult_82_ab_8__33_, u5_mult_82_ab_8__34_,
         u5_mult_82_ab_8__35_, u5_mult_82_ab_8__36_, u5_mult_82_ab_8__37_,
         u5_mult_82_ab_8__38_, u5_mult_82_ab_8__39_, u5_mult_82_ab_8__40_,
         u5_mult_82_ab_8__41_, u5_mult_82_ab_8__42_, u5_mult_82_ab_8__43_,
         u5_mult_82_ab_8__44_, u5_mult_82_ab_8__45_, u5_mult_82_ab_8__46_,
         u5_mult_82_ab_8__47_, u5_mult_82_ab_8__48_, u5_mult_82_ab_8__49_,
         u5_mult_82_ab_8__50_, u5_mult_82_ab_8__51_, u5_mult_82_ab_8__52_,
         u5_mult_82_ab_9__0_, u5_mult_82_ab_9__1_, u5_mult_82_ab_9__2_,
         u5_mult_82_ab_9__3_, u5_mult_82_ab_9__4_, u5_mult_82_ab_9__5_,
         u5_mult_82_ab_9__6_, u5_mult_82_ab_9__7_, u5_mult_82_ab_9__8_,
         u5_mult_82_ab_9__9_, u5_mult_82_ab_9__10_, u5_mult_82_ab_9__11_,
         u5_mult_82_ab_9__12_, u5_mult_82_ab_9__13_, u5_mult_82_ab_9__14_,
         u5_mult_82_ab_9__15_, u5_mult_82_ab_9__16_, u5_mult_82_ab_9__17_,
         u5_mult_82_ab_9__18_, u5_mult_82_ab_9__19_, u5_mult_82_ab_9__20_,
         u5_mult_82_ab_9__21_, u5_mult_82_ab_9__22_, u5_mult_82_ab_9__23_,
         u5_mult_82_ab_9__24_, u5_mult_82_ab_9__25_, u5_mult_82_ab_9__26_,
         u5_mult_82_ab_9__27_, u5_mult_82_ab_9__28_, u5_mult_82_ab_9__29_,
         u5_mult_82_ab_9__30_, u5_mult_82_ab_9__31_, u5_mult_82_ab_9__32_,
         u5_mult_82_ab_9__33_, u5_mult_82_ab_9__34_, u5_mult_82_ab_9__35_,
         u5_mult_82_ab_9__36_, u5_mult_82_ab_9__37_, u5_mult_82_ab_9__38_,
         u5_mult_82_ab_9__39_, u5_mult_82_ab_9__40_, u5_mult_82_ab_9__41_,
         u5_mult_82_ab_9__42_, u5_mult_82_ab_9__43_, u5_mult_82_ab_9__44_,
         u5_mult_82_ab_9__45_, u5_mult_82_ab_9__46_, u5_mult_82_ab_9__47_,
         u5_mult_82_ab_9__48_, u5_mult_82_ab_9__49_, u5_mult_82_ab_9__50_,
         u5_mult_82_ab_9__51_, u5_mult_82_ab_9__52_, u5_mult_82_ab_10__0_,
         u5_mult_82_ab_10__1_, u5_mult_82_ab_10__2_, u5_mult_82_ab_10__3_,
         u5_mult_82_ab_10__4_, u5_mult_82_ab_10__5_, u5_mult_82_ab_10__6_,
         u5_mult_82_ab_10__7_, u5_mult_82_ab_10__8_, u5_mult_82_ab_10__9_,
         u5_mult_82_ab_10__10_, u5_mult_82_ab_10__11_, u5_mult_82_ab_10__12_,
         u5_mult_82_ab_10__13_, u5_mult_82_ab_10__14_, u5_mult_82_ab_10__15_,
         u5_mult_82_ab_10__16_, u5_mult_82_ab_10__17_, u5_mult_82_ab_10__18_,
         u5_mult_82_ab_10__19_, u5_mult_82_ab_10__20_, u5_mult_82_ab_10__21_,
         u5_mult_82_ab_10__22_, u5_mult_82_ab_10__23_, u5_mult_82_ab_10__24_,
         u5_mult_82_ab_10__25_, u5_mult_82_ab_10__26_, u5_mult_82_ab_10__27_,
         u5_mult_82_ab_10__28_, u5_mult_82_ab_10__29_, u5_mult_82_ab_10__30_,
         u5_mult_82_ab_10__31_, u5_mult_82_ab_10__32_, u5_mult_82_ab_10__33_,
         u5_mult_82_ab_10__34_, u5_mult_82_ab_10__35_, u5_mult_82_ab_10__36_,
         u5_mult_82_ab_10__37_, u5_mult_82_ab_10__38_, u5_mult_82_ab_10__39_,
         u5_mult_82_ab_10__40_, u5_mult_82_ab_10__41_, u5_mult_82_ab_10__42_,
         u5_mult_82_ab_10__43_, u5_mult_82_ab_10__44_, u5_mult_82_ab_10__45_,
         u5_mult_82_ab_10__46_, u5_mult_82_ab_10__47_, u5_mult_82_ab_10__48_,
         u5_mult_82_ab_10__49_, u5_mult_82_ab_10__50_, u5_mult_82_ab_10__51_,
         u5_mult_82_ab_10__52_, u5_mult_82_ab_11__0_, u5_mult_82_ab_11__1_,
         u5_mult_82_ab_11__2_, u5_mult_82_ab_11__3_, u5_mult_82_ab_11__4_,
         u5_mult_82_ab_11__5_, u5_mult_82_ab_11__6_, u5_mult_82_ab_11__7_,
         u5_mult_82_ab_11__8_, u5_mult_82_ab_11__9_, u5_mult_82_ab_11__10_,
         u5_mult_82_ab_11__11_, u5_mult_82_ab_11__12_, u5_mult_82_ab_11__13_,
         u5_mult_82_ab_11__14_, u5_mult_82_ab_11__15_, u5_mult_82_ab_11__16_,
         u5_mult_82_ab_11__17_, u5_mult_82_ab_11__18_, u5_mult_82_ab_11__19_,
         u5_mult_82_ab_11__20_, u5_mult_82_ab_11__21_, u5_mult_82_ab_11__22_,
         u5_mult_82_ab_11__23_, u5_mult_82_ab_11__24_, u5_mult_82_ab_11__25_,
         u5_mult_82_ab_11__26_, u5_mult_82_ab_11__27_, u5_mult_82_ab_11__28_,
         u5_mult_82_ab_11__29_, u5_mult_82_ab_11__30_, u5_mult_82_ab_11__31_,
         u5_mult_82_ab_11__32_, u5_mult_82_ab_11__33_, u5_mult_82_ab_11__34_,
         u5_mult_82_ab_11__35_, u5_mult_82_ab_11__36_, u5_mult_82_ab_11__37_,
         u5_mult_82_ab_11__38_, u5_mult_82_ab_11__39_, u5_mult_82_ab_11__40_,
         u5_mult_82_ab_11__41_, u5_mult_82_ab_11__42_, u5_mult_82_ab_11__43_,
         u5_mult_82_ab_11__44_, u5_mult_82_ab_11__45_, u5_mult_82_ab_11__46_,
         u5_mult_82_ab_11__47_, u5_mult_82_ab_11__48_, u5_mult_82_ab_11__49_,
         u5_mult_82_ab_11__50_, u5_mult_82_ab_11__51_, u5_mult_82_ab_11__52_,
         u5_mult_82_ab_12__0_, u5_mult_82_ab_12__1_, u5_mult_82_ab_12__2_,
         u5_mult_82_ab_12__3_, u5_mult_82_ab_12__4_, u5_mult_82_ab_12__5_,
         u5_mult_82_ab_12__6_, u5_mult_82_ab_12__7_, u5_mult_82_ab_12__8_,
         u5_mult_82_ab_12__9_, u5_mult_82_ab_12__10_, u5_mult_82_ab_12__11_,
         u5_mult_82_ab_12__12_, u5_mult_82_ab_12__13_, u5_mult_82_ab_12__14_,
         u5_mult_82_ab_12__15_, u5_mult_82_ab_12__16_, u5_mult_82_ab_12__17_,
         u5_mult_82_ab_12__18_, u5_mult_82_ab_12__19_, u5_mult_82_ab_12__20_,
         u5_mult_82_ab_12__21_, u5_mult_82_ab_12__22_, u5_mult_82_ab_12__23_,
         u5_mult_82_ab_12__24_, u5_mult_82_ab_12__25_, u5_mult_82_ab_12__26_,
         u5_mult_82_ab_12__27_, u5_mult_82_ab_12__28_, u5_mult_82_ab_12__29_,
         u5_mult_82_ab_12__30_, u5_mult_82_ab_12__31_, u5_mult_82_ab_12__32_,
         u5_mult_82_ab_12__33_, u5_mult_82_ab_12__34_, u5_mult_82_ab_12__35_,
         u5_mult_82_ab_12__36_, u5_mult_82_ab_12__37_, u5_mult_82_ab_12__38_,
         u5_mult_82_ab_12__39_, u5_mult_82_ab_12__40_, u5_mult_82_ab_12__41_,
         u5_mult_82_ab_12__42_, u5_mult_82_ab_12__43_, u5_mult_82_ab_12__44_,
         u5_mult_82_ab_12__45_, u5_mult_82_ab_12__46_, u5_mult_82_ab_12__47_,
         u5_mult_82_ab_12__48_, u5_mult_82_ab_12__49_, u5_mult_82_ab_12__50_,
         u5_mult_82_ab_12__51_, u5_mult_82_ab_12__52_, u5_mult_82_ab_13__0_,
         u5_mult_82_ab_13__1_, u5_mult_82_ab_13__2_, u5_mult_82_ab_13__3_,
         u5_mult_82_ab_13__4_, u5_mult_82_ab_13__5_, u5_mult_82_ab_13__6_,
         u5_mult_82_ab_13__7_, u5_mult_82_ab_13__8_, u5_mult_82_ab_13__9_,
         u5_mult_82_ab_13__10_, u5_mult_82_ab_13__11_, u5_mult_82_ab_13__12_,
         u5_mult_82_ab_13__13_, u5_mult_82_ab_13__14_, u5_mult_82_ab_13__15_,
         u5_mult_82_ab_13__16_, u5_mult_82_ab_13__17_, u5_mult_82_ab_13__18_,
         u5_mult_82_ab_13__19_, u5_mult_82_ab_13__20_, u5_mult_82_ab_13__21_,
         u5_mult_82_ab_13__22_, u5_mult_82_ab_13__23_, u5_mult_82_ab_13__24_,
         u5_mult_82_ab_13__25_, u5_mult_82_ab_13__26_, u5_mult_82_ab_13__27_,
         u5_mult_82_ab_13__28_, u5_mult_82_ab_13__29_, u5_mult_82_ab_13__30_,
         u5_mult_82_ab_13__31_, u5_mult_82_ab_13__32_, u5_mult_82_ab_13__33_,
         u5_mult_82_ab_13__34_, u5_mult_82_ab_13__35_, u5_mult_82_ab_13__36_,
         u5_mult_82_ab_13__37_, u5_mult_82_ab_13__38_, u5_mult_82_ab_13__39_,
         u5_mult_82_ab_13__40_, u5_mult_82_ab_13__41_, u5_mult_82_ab_13__42_,
         u5_mult_82_ab_13__43_, u5_mult_82_ab_13__44_, u5_mult_82_ab_13__45_,
         u5_mult_82_ab_13__46_, u5_mult_82_ab_13__47_, u5_mult_82_ab_13__48_,
         u5_mult_82_ab_13__49_, u5_mult_82_ab_13__50_, u5_mult_82_ab_13__51_,
         u5_mult_82_ab_13__52_, u5_mult_82_ab_14__0_, u5_mult_82_ab_14__1_,
         u5_mult_82_ab_14__2_, u5_mult_82_ab_14__3_, u5_mult_82_ab_14__4_,
         u5_mult_82_ab_14__5_, u5_mult_82_ab_14__6_, u5_mult_82_ab_14__7_,
         u5_mult_82_ab_14__8_, u5_mult_82_ab_14__9_, u5_mult_82_ab_14__10_,
         u5_mult_82_ab_14__11_, u5_mult_82_ab_14__12_, u5_mult_82_ab_14__13_,
         u5_mult_82_ab_14__14_, u5_mult_82_ab_14__15_, u5_mult_82_ab_14__16_,
         u5_mult_82_ab_14__17_, u5_mult_82_ab_14__18_, u5_mult_82_ab_14__19_,
         u5_mult_82_ab_14__20_, u5_mult_82_ab_14__21_, u5_mult_82_ab_14__22_,
         u5_mult_82_ab_14__23_, u5_mult_82_ab_14__24_, u5_mult_82_ab_14__25_,
         u5_mult_82_ab_14__26_, u5_mult_82_ab_14__27_, u5_mult_82_ab_14__28_,
         u5_mult_82_ab_14__29_, u5_mult_82_ab_14__30_, u5_mult_82_ab_14__31_,
         u5_mult_82_ab_14__32_, u5_mult_82_ab_14__33_, u5_mult_82_ab_14__34_,
         u5_mult_82_ab_14__35_, u5_mult_82_ab_14__36_, u5_mult_82_ab_14__37_,
         u5_mult_82_ab_14__38_, u5_mult_82_ab_14__39_, u5_mult_82_ab_14__40_,
         u5_mult_82_ab_14__41_, u5_mult_82_ab_14__42_, u5_mult_82_ab_14__43_,
         u5_mult_82_ab_14__44_, u5_mult_82_ab_14__45_, u5_mult_82_ab_14__46_,
         u5_mult_82_ab_14__47_, u5_mult_82_ab_14__48_, u5_mult_82_ab_14__49_,
         u5_mult_82_ab_14__50_, u5_mult_82_ab_14__51_, u5_mult_82_ab_14__52_,
         u5_mult_82_ab_15__0_, u5_mult_82_ab_15__1_, u5_mult_82_ab_15__2_,
         u5_mult_82_ab_15__3_, u5_mult_82_ab_15__4_, u5_mult_82_ab_15__5_,
         u5_mult_82_ab_15__6_, u5_mult_82_ab_15__7_, u5_mult_82_ab_15__8_,
         u5_mult_82_ab_15__9_, u5_mult_82_ab_15__10_, u5_mult_82_ab_15__11_,
         u5_mult_82_ab_15__12_, u5_mult_82_ab_15__13_, u5_mult_82_ab_15__14_,
         u5_mult_82_ab_15__15_, u5_mult_82_ab_15__16_, u5_mult_82_ab_15__17_,
         u5_mult_82_ab_15__18_, u5_mult_82_ab_15__19_, u5_mult_82_ab_15__20_,
         u5_mult_82_ab_15__21_, u5_mult_82_ab_15__22_, u5_mult_82_ab_15__23_,
         u5_mult_82_ab_15__24_, u5_mult_82_ab_15__25_, u5_mult_82_ab_15__26_,
         u5_mult_82_ab_15__27_, u5_mult_82_ab_15__28_, u5_mult_82_ab_15__29_,
         u5_mult_82_ab_15__30_, u5_mult_82_ab_15__31_, u5_mult_82_ab_15__32_,
         u5_mult_82_ab_15__33_, u5_mult_82_ab_15__34_, u5_mult_82_ab_15__35_,
         u5_mult_82_ab_15__36_, u5_mult_82_ab_15__37_, u5_mult_82_ab_15__38_,
         u5_mult_82_ab_15__39_, u5_mult_82_ab_15__40_, u5_mult_82_ab_15__41_,
         u5_mult_82_ab_15__42_, u5_mult_82_ab_15__43_, u5_mult_82_ab_15__44_,
         u5_mult_82_ab_15__45_, u5_mult_82_ab_15__46_, u5_mult_82_ab_15__47_,
         u5_mult_82_ab_15__48_, u5_mult_82_ab_15__49_, u5_mult_82_ab_15__50_,
         u5_mult_82_ab_15__51_, u5_mult_82_ab_15__52_, u5_mult_82_ab_16__0_,
         u5_mult_82_ab_16__1_, u5_mult_82_ab_16__2_, u5_mult_82_ab_16__3_,
         u5_mult_82_ab_16__4_, u5_mult_82_ab_16__5_, u5_mult_82_ab_16__6_,
         u5_mult_82_ab_16__7_, u5_mult_82_ab_16__8_, u5_mult_82_ab_16__9_,
         u5_mult_82_ab_16__10_, u5_mult_82_ab_16__11_, u5_mult_82_ab_16__12_,
         u5_mult_82_ab_16__13_, u5_mult_82_ab_16__14_, u5_mult_82_ab_16__15_,
         u5_mult_82_ab_16__16_, u5_mult_82_ab_16__17_, u5_mult_82_ab_16__18_,
         u5_mult_82_ab_16__19_, u5_mult_82_ab_16__20_, u5_mult_82_ab_16__21_,
         u5_mult_82_ab_16__22_, u5_mult_82_ab_16__23_, u5_mult_82_ab_16__24_,
         u5_mult_82_ab_16__25_, u5_mult_82_ab_16__26_, u5_mult_82_ab_16__27_,
         u5_mult_82_ab_16__28_, u5_mult_82_ab_16__29_, u5_mult_82_ab_16__30_,
         u5_mult_82_ab_16__31_, u5_mult_82_ab_16__32_, u5_mult_82_ab_16__33_,
         u5_mult_82_ab_16__34_, u5_mult_82_ab_16__35_, u5_mult_82_ab_16__36_,
         u5_mult_82_ab_16__37_, u5_mult_82_ab_16__38_, u5_mult_82_ab_16__39_,
         u5_mult_82_ab_16__40_, u5_mult_82_ab_16__41_, u5_mult_82_ab_16__42_,
         u5_mult_82_ab_16__43_, u5_mult_82_ab_16__44_, u5_mult_82_ab_16__45_,
         u5_mult_82_ab_16__46_, u5_mult_82_ab_16__47_, u5_mult_82_ab_16__48_,
         u5_mult_82_ab_16__49_, u5_mult_82_ab_16__50_, u5_mult_82_ab_16__51_,
         u5_mult_82_ab_16__52_, u5_mult_82_ab_17__0_, u5_mult_82_ab_17__1_,
         u5_mult_82_ab_17__2_, u5_mult_82_ab_17__3_, u5_mult_82_ab_17__4_,
         u5_mult_82_ab_17__5_, u5_mult_82_ab_17__6_, u5_mult_82_ab_17__7_,
         u5_mult_82_ab_17__8_, u5_mult_82_ab_17__9_, u5_mult_82_ab_17__10_,
         u5_mult_82_ab_17__11_, u5_mult_82_ab_17__12_, u5_mult_82_ab_17__13_,
         u5_mult_82_ab_17__14_, u5_mult_82_ab_17__15_, u5_mult_82_ab_17__16_,
         u5_mult_82_ab_17__17_, u5_mult_82_ab_17__18_, u5_mult_82_ab_17__19_,
         u5_mult_82_ab_17__20_, u5_mult_82_ab_17__21_, u5_mult_82_ab_17__22_,
         u5_mult_82_ab_17__23_, u5_mult_82_ab_17__24_, u5_mult_82_ab_17__25_,
         u5_mult_82_ab_17__26_, u5_mult_82_ab_17__27_, u5_mult_82_ab_17__28_,
         u5_mult_82_ab_17__29_, u5_mult_82_ab_17__30_, u5_mult_82_ab_17__31_,
         u5_mult_82_ab_17__32_, u5_mult_82_ab_17__33_, u5_mult_82_ab_17__34_,
         u5_mult_82_ab_17__35_, u5_mult_82_ab_17__36_, u5_mult_82_ab_17__37_,
         u5_mult_82_ab_17__38_, u5_mult_82_ab_17__39_, u5_mult_82_ab_17__40_,
         u5_mult_82_ab_17__41_, u5_mult_82_ab_17__42_, u5_mult_82_ab_17__43_,
         u5_mult_82_ab_17__44_, u5_mult_82_ab_17__45_, u5_mult_82_ab_17__46_,
         u5_mult_82_ab_17__47_, u5_mult_82_ab_17__48_, u5_mult_82_ab_17__49_,
         u5_mult_82_ab_17__50_, u5_mult_82_ab_17__51_, u5_mult_82_ab_17__52_,
         u5_mult_82_ab_18__0_, u5_mult_82_ab_18__1_, u5_mult_82_ab_18__2_,
         u5_mult_82_ab_18__3_, u5_mult_82_ab_18__4_, u5_mult_82_ab_18__5_,
         u5_mult_82_ab_18__6_, u5_mult_82_ab_18__7_, u5_mult_82_ab_18__8_,
         u5_mult_82_ab_18__9_, u5_mult_82_ab_18__10_, u5_mult_82_ab_18__11_,
         u5_mult_82_ab_18__12_, u5_mult_82_ab_18__13_, u5_mult_82_ab_18__14_,
         u5_mult_82_ab_18__15_, u5_mult_82_ab_18__16_, u5_mult_82_ab_18__17_,
         u5_mult_82_ab_18__18_, u5_mult_82_ab_18__19_, u5_mult_82_ab_18__20_,
         u5_mult_82_ab_18__21_, u5_mult_82_ab_18__22_, u5_mult_82_ab_18__23_,
         u5_mult_82_ab_18__24_, u5_mult_82_ab_18__25_, u5_mult_82_ab_18__26_,
         u5_mult_82_ab_18__27_, u5_mult_82_ab_18__28_, u5_mult_82_ab_18__29_,
         u5_mult_82_ab_18__30_, u5_mult_82_ab_18__31_, u5_mult_82_ab_18__32_,
         u5_mult_82_ab_18__33_, u5_mult_82_ab_18__34_, u5_mult_82_ab_18__35_,
         u5_mult_82_ab_18__36_, u5_mult_82_ab_18__37_, u5_mult_82_ab_18__38_,
         u5_mult_82_ab_18__39_, u5_mult_82_ab_18__40_, u5_mult_82_ab_18__41_,
         u5_mult_82_ab_18__42_, u5_mult_82_ab_18__43_, u5_mult_82_ab_18__44_,
         u5_mult_82_ab_18__45_, u5_mult_82_ab_18__46_, u5_mult_82_ab_18__47_,
         u5_mult_82_ab_18__48_, u5_mult_82_ab_18__49_, u5_mult_82_ab_18__50_,
         u5_mult_82_ab_18__51_, u5_mult_82_ab_18__52_, u5_mult_82_ab_19__0_,
         u5_mult_82_ab_19__1_, u5_mult_82_ab_19__2_, u5_mult_82_ab_19__3_,
         u5_mult_82_ab_19__4_, u5_mult_82_ab_19__5_, u5_mult_82_ab_19__6_,
         u5_mult_82_ab_19__7_, u5_mult_82_ab_19__8_, u5_mult_82_ab_19__9_,
         u5_mult_82_ab_19__10_, u5_mult_82_ab_19__11_, u5_mult_82_ab_19__12_,
         u5_mult_82_ab_19__13_, u5_mult_82_ab_19__14_, u5_mult_82_ab_19__15_,
         u5_mult_82_ab_19__16_, u5_mult_82_ab_19__17_, u5_mult_82_ab_19__18_,
         u5_mult_82_ab_19__19_, u5_mult_82_ab_19__20_, u5_mult_82_ab_19__21_,
         u5_mult_82_ab_19__22_, u5_mult_82_ab_19__23_, u5_mult_82_ab_19__24_,
         u5_mult_82_ab_19__25_, u5_mult_82_ab_19__26_, u5_mult_82_ab_19__27_,
         u5_mult_82_ab_19__28_, u5_mult_82_ab_19__29_, u5_mult_82_ab_19__30_,
         u5_mult_82_ab_19__31_, u5_mult_82_ab_19__32_, u5_mult_82_ab_19__33_,
         u5_mult_82_ab_19__34_, u5_mult_82_ab_19__35_, u5_mult_82_ab_19__36_,
         u5_mult_82_ab_19__37_, u5_mult_82_ab_19__38_, u5_mult_82_ab_19__39_,
         u5_mult_82_ab_19__40_, u5_mult_82_ab_19__41_, u5_mult_82_ab_19__42_,
         u5_mult_82_ab_19__43_, u5_mult_82_ab_19__44_, u5_mult_82_ab_19__45_,
         u5_mult_82_ab_19__46_, u5_mult_82_ab_19__47_, u5_mult_82_ab_19__48_,
         u5_mult_82_ab_19__49_, u5_mult_82_ab_19__50_, u5_mult_82_ab_19__51_,
         u5_mult_82_ab_19__52_, u5_mult_82_ab_20__0_, u5_mult_82_ab_20__1_,
         u5_mult_82_ab_20__2_, u5_mult_82_ab_20__3_, u5_mult_82_ab_20__4_,
         u5_mult_82_ab_20__5_, u5_mult_82_ab_20__6_, u5_mult_82_ab_20__7_,
         u5_mult_82_ab_20__8_, u5_mult_82_ab_20__9_, u5_mult_82_ab_20__10_,
         u5_mult_82_ab_20__11_, u5_mult_82_ab_20__12_, u5_mult_82_ab_20__13_,
         u5_mult_82_ab_20__14_, u5_mult_82_ab_20__15_, u5_mult_82_ab_20__16_,
         u5_mult_82_ab_20__17_, u5_mult_82_ab_20__18_, u5_mult_82_ab_20__19_,
         u5_mult_82_ab_20__20_, u5_mult_82_ab_20__21_, u5_mult_82_ab_20__22_,
         u5_mult_82_ab_20__23_, u5_mult_82_ab_20__24_, u5_mult_82_ab_20__25_,
         u5_mult_82_ab_20__26_, u5_mult_82_ab_20__27_, u5_mult_82_ab_20__28_,
         u5_mult_82_ab_20__29_, u5_mult_82_ab_20__30_, u5_mult_82_ab_20__31_,
         u5_mult_82_ab_20__32_, u5_mult_82_ab_20__33_, u5_mult_82_ab_20__34_,
         u5_mult_82_ab_20__35_, u5_mult_82_ab_20__36_, u5_mult_82_ab_20__37_,
         u5_mult_82_ab_20__38_, u5_mult_82_ab_20__39_, u5_mult_82_ab_20__40_,
         u5_mult_82_ab_20__41_, u5_mult_82_ab_20__42_, u5_mult_82_ab_20__43_,
         u5_mult_82_ab_20__44_, u5_mult_82_ab_20__45_, u5_mult_82_ab_20__46_,
         u5_mult_82_ab_20__47_, u5_mult_82_ab_20__48_, u5_mult_82_ab_20__49_,
         u5_mult_82_ab_20__50_, u5_mult_82_ab_20__51_, u5_mult_82_ab_20__52_,
         u5_mult_82_ab_21__0_, u5_mult_82_ab_21__1_, u5_mult_82_ab_21__2_,
         u5_mult_82_ab_21__3_, u5_mult_82_ab_21__4_, u5_mult_82_ab_21__5_,
         u5_mult_82_ab_21__6_, u5_mult_82_ab_21__7_, u5_mult_82_ab_21__8_,
         u5_mult_82_ab_21__9_, u5_mult_82_ab_21__10_, u5_mult_82_ab_21__11_,
         u5_mult_82_ab_21__12_, u5_mult_82_ab_21__13_, u5_mult_82_ab_21__14_,
         u5_mult_82_ab_21__15_, u5_mult_82_ab_21__16_, u5_mult_82_ab_21__17_,
         u5_mult_82_ab_21__18_, u5_mult_82_ab_21__19_, u5_mult_82_ab_21__20_,
         u5_mult_82_ab_21__21_, u5_mult_82_ab_21__22_, u5_mult_82_ab_21__23_,
         u5_mult_82_ab_21__24_, u5_mult_82_ab_21__25_, u5_mult_82_ab_21__26_,
         u5_mult_82_ab_21__27_, u5_mult_82_ab_21__28_, u5_mult_82_ab_21__29_,
         u5_mult_82_ab_21__30_, u5_mult_82_ab_21__31_, u5_mult_82_ab_21__32_,
         u5_mult_82_ab_21__33_, u5_mult_82_ab_21__34_, u5_mult_82_ab_21__35_,
         u5_mult_82_ab_21__36_, u5_mult_82_ab_21__37_, u5_mult_82_ab_21__38_,
         u5_mult_82_ab_21__39_, u5_mult_82_ab_21__40_, u5_mult_82_ab_21__41_,
         u5_mult_82_ab_21__42_, u5_mult_82_ab_21__43_, u5_mult_82_ab_21__44_,
         u5_mult_82_ab_21__45_, u5_mult_82_ab_21__46_, u5_mult_82_ab_21__47_,
         u5_mult_82_ab_21__48_, u5_mult_82_ab_21__49_, u5_mult_82_ab_21__50_,
         u5_mult_82_ab_21__51_, u5_mult_82_ab_21__52_, u5_mult_82_ab_22__0_,
         u5_mult_82_ab_22__1_, u5_mult_82_ab_22__2_, u5_mult_82_ab_22__3_,
         u5_mult_82_ab_22__4_, u5_mult_82_ab_22__5_, u5_mult_82_ab_22__6_,
         u5_mult_82_ab_22__7_, u5_mult_82_ab_22__8_, u5_mult_82_ab_22__9_,
         u5_mult_82_ab_22__10_, u5_mult_82_ab_22__11_, u5_mult_82_ab_22__12_,
         u5_mult_82_ab_22__13_, u5_mult_82_ab_22__14_, u5_mult_82_ab_22__15_,
         u5_mult_82_ab_22__16_, u5_mult_82_ab_22__17_, u5_mult_82_ab_22__18_,
         u5_mult_82_ab_22__19_, u5_mult_82_ab_22__20_, u5_mult_82_ab_22__21_,
         u5_mult_82_ab_22__22_, u5_mult_82_ab_22__23_, u5_mult_82_ab_22__24_,
         u5_mult_82_ab_22__25_, u5_mult_82_ab_22__26_, u5_mult_82_ab_22__27_,
         u5_mult_82_ab_22__28_, u5_mult_82_ab_22__29_, u5_mult_82_ab_22__30_,
         u5_mult_82_ab_22__31_, u5_mult_82_ab_22__32_, u5_mult_82_ab_22__33_,
         u5_mult_82_ab_22__34_, u5_mult_82_ab_22__35_, u5_mult_82_ab_22__36_,
         u5_mult_82_ab_22__37_, u5_mult_82_ab_22__38_, u5_mult_82_ab_22__39_,
         u5_mult_82_ab_22__40_, u5_mult_82_ab_22__41_, u5_mult_82_ab_22__42_,
         u5_mult_82_ab_22__43_, u5_mult_82_ab_22__44_, u5_mult_82_ab_22__45_,
         u5_mult_82_ab_22__46_, u5_mult_82_ab_22__47_, u5_mult_82_ab_22__48_,
         u5_mult_82_ab_22__49_, u5_mult_82_ab_22__50_, u5_mult_82_ab_22__51_,
         u5_mult_82_ab_22__52_, u5_mult_82_ab_23__0_, u5_mult_82_ab_23__1_,
         u5_mult_82_ab_23__2_, u5_mult_82_ab_23__3_, u5_mult_82_ab_23__4_,
         u5_mult_82_ab_23__5_, u5_mult_82_ab_23__6_, u5_mult_82_ab_23__7_,
         u5_mult_82_ab_23__8_, u5_mult_82_ab_23__9_, u5_mult_82_ab_23__10_,
         u5_mult_82_ab_23__11_, u5_mult_82_ab_23__12_, u5_mult_82_ab_23__13_,
         u5_mult_82_ab_23__14_, u5_mult_82_ab_23__15_, u5_mult_82_ab_23__16_,
         u5_mult_82_ab_23__17_, u5_mult_82_ab_23__18_, u5_mult_82_ab_23__19_,
         u5_mult_82_ab_23__20_, u5_mult_82_ab_23__21_, u5_mult_82_ab_23__22_,
         u5_mult_82_ab_23__23_, u5_mult_82_ab_23__24_, u5_mult_82_ab_23__25_,
         u5_mult_82_ab_23__26_, u5_mult_82_ab_23__27_, u5_mult_82_ab_23__28_,
         u5_mult_82_ab_23__29_, u5_mult_82_ab_23__30_, u5_mult_82_ab_23__31_,
         u5_mult_82_ab_23__32_, u5_mult_82_ab_23__33_, u5_mult_82_ab_23__34_,
         u5_mult_82_ab_23__35_, u5_mult_82_ab_23__36_, u5_mult_82_ab_23__37_,
         u5_mult_82_ab_23__38_, u5_mult_82_ab_23__39_, u5_mult_82_ab_23__40_,
         u5_mult_82_ab_23__41_, u5_mult_82_ab_23__42_, u5_mult_82_ab_23__43_,
         u5_mult_82_ab_23__44_, u5_mult_82_ab_23__45_, u5_mult_82_ab_23__46_,
         u5_mult_82_ab_23__47_, u5_mult_82_ab_23__48_, u5_mult_82_ab_23__49_,
         u5_mult_82_ab_23__50_, u5_mult_82_ab_23__51_, u5_mult_82_ab_23__52_,
         u5_mult_82_ab_24__0_, u5_mult_82_ab_24__1_, u5_mult_82_ab_24__2_,
         u5_mult_82_ab_24__3_, u5_mult_82_ab_24__4_, u5_mult_82_ab_24__5_,
         u5_mult_82_ab_24__6_, u5_mult_82_ab_24__7_, u5_mult_82_ab_24__8_,
         u5_mult_82_ab_24__9_, u5_mult_82_ab_24__10_, u5_mult_82_ab_24__11_,
         u5_mult_82_ab_24__12_, u5_mult_82_ab_24__13_, u5_mult_82_ab_24__14_,
         u5_mult_82_ab_24__15_, u5_mult_82_ab_24__16_, u5_mult_82_ab_24__17_,
         u5_mult_82_ab_24__18_, u5_mult_82_ab_24__19_, u5_mult_82_ab_24__20_,
         u5_mult_82_ab_24__21_, u5_mult_82_ab_24__22_, u5_mult_82_ab_24__23_,
         u5_mult_82_ab_24__24_, u5_mult_82_ab_24__25_, u5_mult_82_ab_24__26_,
         u5_mult_82_ab_24__27_, u5_mult_82_ab_24__28_, u5_mult_82_ab_24__29_,
         u5_mult_82_ab_24__30_, u5_mult_82_ab_24__31_, u5_mult_82_ab_24__32_,
         u5_mult_82_ab_24__33_, u5_mult_82_ab_24__34_, u5_mult_82_ab_24__35_,
         u5_mult_82_ab_24__36_, u5_mult_82_ab_24__37_, u5_mult_82_ab_24__38_,
         u5_mult_82_ab_24__39_, u5_mult_82_ab_24__40_, u5_mult_82_ab_24__41_,
         u5_mult_82_ab_24__42_, u5_mult_82_ab_24__43_, u5_mult_82_ab_24__44_,
         u5_mult_82_ab_24__45_, u5_mult_82_ab_24__46_, u5_mult_82_ab_24__47_,
         u5_mult_82_ab_24__48_, u5_mult_82_ab_24__49_, u5_mult_82_ab_24__50_,
         u5_mult_82_ab_24__51_, u5_mult_82_ab_24__52_, u5_mult_82_ab_25__0_,
         u5_mult_82_ab_25__1_, u5_mult_82_ab_25__2_, u5_mult_82_ab_25__3_,
         u5_mult_82_ab_25__4_, u5_mult_82_ab_25__5_, u5_mult_82_ab_25__6_,
         u5_mult_82_ab_25__7_, u5_mult_82_ab_25__8_, u5_mult_82_ab_25__9_,
         u5_mult_82_ab_25__10_, u5_mult_82_ab_25__11_, u5_mult_82_ab_25__12_,
         u5_mult_82_ab_25__13_, u5_mult_82_ab_25__14_, u5_mult_82_ab_25__15_,
         u5_mult_82_ab_25__16_, u5_mult_82_ab_25__17_, u5_mult_82_ab_25__18_,
         u5_mult_82_ab_25__19_, u5_mult_82_ab_25__20_, u5_mult_82_ab_25__21_,
         u5_mult_82_ab_25__22_, u5_mult_82_ab_25__23_, u5_mult_82_ab_25__24_,
         u5_mult_82_ab_25__25_, u5_mult_82_ab_25__26_, u5_mult_82_ab_25__27_,
         u5_mult_82_ab_25__28_, u5_mult_82_ab_25__29_, u5_mult_82_ab_25__30_,
         u5_mult_82_ab_25__31_, u5_mult_82_ab_25__32_, u5_mult_82_ab_25__33_,
         u5_mult_82_ab_25__34_, u5_mult_82_ab_25__35_, u5_mult_82_ab_25__36_,
         u5_mult_82_ab_25__37_, u5_mult_82_ab_25__38_, u5_mult_82_ab_25__39_,
         u5_mult_82_ab_25__40_, u5_mult_82_ab_25__41_, u5_mult_82_ab_25__42_,
         u5_mult_82_ab_25__43_, u5_mult_82_ab_25__44_, u5_mult_82_ab_25__45_,
         u5_mult_82_ab_25__46_, u5_mult_82_ab_25__47_, u5_mult_82_ab_25__48_,
         u5_mult_82_ab_25__49_, u5_mult_82_ab_25__50_, u5_mult_82_ab_25__51_,
         u5_mult_82_ab_25__52_, u5_mult_82_ab_26__0_, u5_mult_82_ab_26__1_,
         u5_mult_82_ab_26__2_, u5_mult_82_ab_26__3_, u5_mult_82_ab_26__4_,
         u5_mult_82_ab_26__5_, u5_mult_82_ab_26__6_, u5_mult_82_ab_26__7_,
         u5_mult_82_ab_26__8_, u5_mult_82_ab_26__9_, u5_mult_82_ab_26__10_,
         u5_mult_82_ab_26__11_, u5_mult_82_ab_26__12_, u5_mult_82_ab_26__13_,
         u5_mult_82_ab_26__14_, u5_mult_82_ab_26__15_, u5_mult_82_ab_26__16_,
         u5_mult_82_ab_26__17_, u5_mult_82_ab_26__18_, u5_mult_82_ab_26__19_,
         u5_mult_82_ab_26__20_, u5_mult_82_ab_26__21_, u5_mult_82_ab_26__22_,
         u5_mult_82_ab_26__23_, u5_mult_82_ab_26__24_, u5_mult_82_ab_26__25_,
         u5_mult_82_ab_26__26_, u5_mult_82_ab_26__27_, u5_mult_82_ab_26__28_,
         u5_mult_82_ab_26__29_, u5_mult_82_ab_26__30_, u5_mult_82_ab_26__31_,
         u5_mult_82_ab_26__32_, u5_mult_82_ab_26__33_, u5_mult_82_ab_26__34_,
         u5_mult_82_ab_26__35_, u5_mult_82_ab_26__36_, u5_mult_82_ab_26__37_,
         u5_mult_82_ab_26__38_, u5_mult_82_ab_26__39_, u5_mult_82_ab_26__40_,
         u5_mult_82_ab_26__41_, u5_mult_82_ab_26__42_, u5_mult_82_ab_26__43_,
         u5_mult_82_ab_26__44_, u5_mult_82_ab_26__45_, u5_mult_82_ab_26__46_,
         u5_mult_82_ab_26__47_, u5_mult_82_ab_26__48_, u5_mult_82_ab_26__49_,
         u5_mult_82_ab_26__50_, u5_mult_82_ab_26__51_, u5_mult_82_ab_26__52_,
         u5_mult_82_ab_27__0_, u5_mult_82_ab_27__1_, u5_mult_82_ab_27__2_,
         u5_mult_82_ab_27__3_, u5_mult_82_ab_27__4_, u5_mult_82_ab_27__5_,
         u5_mult_82_ab_27__6_, u5_mult_82_ab_27__7_, u5_mult_82_ab_27__8_,
         u5_mult_82_ab_27__9_, u5_mult_82_ab_27__10_, u5_mult_82_ab_27__11_,
         u5_mult_82_ab_27__12_, u5_mult_82_ab_27__13_, u5_mult_82_ab_27__14_,
         u5_mult_82_ab_27__15_, u5_mult_82_ab_27__16_, u5_mult_82_ab_27__17_,
         u5_mult_82_ab_27__18_, u5_mult_82_ab_27__19_, u5_mult_82_ab_27__20_,
         u5_mult_82_ab_27__21_, u5_mult_82_ab_27__22_, u5_mult_82_ab_27__23_,
         u5_mult_82_ab_27__24_, u5_mult_82_ab_27__25_, u5_mult_82_ab_27__26_,
         u5_mult_82_ab_27__27_, u5_mult_82_ab_27__28_, u5_mult_82_ab_27__29_,
         u5_mult_82_ab_27__30_, u5_mult_82_ab_27__31_, u5_mult_82_ab_27__32_,
         u5_mult_82_ab_27__33_, u5_mult_82_ab_27__34_, u5_mult_82_ab_27__35_,
         u5_mult_82_ab_27__36_, u5_mult_82_ab_27__37_, u5_mult_82_ab_27__38_,
         u5_mult_82_ab_27__39_, u5_mult_82_ab_27__40_, u5_mult_82_ab_27__41_,
         u5_mult_82_ab_27__42_, u5_mult_82_ab_27__43_, u5_mult_82_ab_27__44_,
         u5_mult_82_ab_27__45_, u5_mult_82_ab_27__46_, u5_mult_82_ab_27__47_,
         u5_mult_82_ab_27__48_, u5_mult_82_ab_27__49_, u5_mult_82_ab_27__50_,
         u5_mult_82_ab_27__51_, u5_mult_82_ab_27__52_, u5_mult_82_ab_28__0_,
         u5_mult_82_ab_28__1_, u5_mult_82_ab_28__2_, u5_mult_82_ab_28__3_,
         u5_mult_82_ab_28__4_, u5_mult_82_ab_28__5_, u5_mult_82_ab_28__6_,
         u5_mult_82_ab_28__7_, u5_mult_82_ab_28__8_, u5_mult_82_ab_28__9_,
         u5_mult_82_ab_28__10_, u5_mult_82_ab_28__11_, u5_mult_82_ab_28__12_,
         u5_mult_82_ab_28__13_, u5_mult_82_ab_28__14_, u5_mult_82_ab_28__15_,
         u5_mult_82_ab_28__16_, u5_mult_82_ab_28__17_, u5_mult_82_ab_28__18_,
         u5_mult_82_ab_28__19_, u5_mult_82_ab_28__20_, u5_mult_82_ab_28__21_,
         u5_mult_82_ab_28__22_, u5_mult_82_ab_28__23_, u5_mult_82_ab_28__24_,
         u5_mult_82_ab_28__25_, u5_mult_82_ab_28__26_, u5_mult_82_ab_28__27_,
         u5_mult_82_ab_28__28_, u5_mult_82_ab_28__29_, u5_mult_82_ab_28__30_,
         u5_mult_82_ab_28__31_, u5_mult_82_ab_28__32_, u5_mult_82_ab_28__33_,
         u5_mult_82_ab_28__34_, u5_mult_82_ab_28__35_, u5_mult_82_ab_28__36_,
         u5_mult_82_ab_28__37_, u5_mult_82_ab_28__38_, u5_mult_82_ab_28__39_,
         u5_mult_82_ab_28__40_, u5_mult_82_ab_28__41_, u5_mult_82_ab_28__42_,
         u5_mult_82_ab_28__43_, u5_mult_82_ab_28__44_, u5_mult_82_ab_28__45_,
         u5_mult_82_ab_28__46_, u5_mult_82_ab_28__47_, u5_mult_82_ab_28__48_,
         u5_mult_82_ab_28__49_, u5_mult_82_ab_28__50_, u5_mult_82_ab_28__51_,
         u5_mult_82_ab_28__52_, u5_mult_82_ab_29__0_, u5_mult_82_ab_29__1_,
         u5_mult_82_ab_29__2_, u5_mult_82_ab_29__3_, u5_mult_82_ab_29__4_,
         u5_mult_82_ab_29__5_, u5_mult_82_ab_29__6_, u5_mult_82_ab_29__7_,
         u5_mult_82_ab_29__8_, u5_mult_82_ab_29__9_, u5_mult_82_ab_29__10_,
         u5_mult_82_ab_29__11_, u5_mult_82_ab_29__12_, u5_mult_82_ab_29__13_,
         u5_mult_82_ab_29__14_, u5_mult_82_ab_29__15_, u5_mult_82_ab_29__16_,
         u5_mult_82_ab_29__17_, u5_mult_82_ab_29__18_, u5_mult_82_ab_29__19_,
         u5_mult_82_ab_29__20_, u5_mult_82_ab_29__21_, u5_mult_82_ab_29__22_,
         u5_mult_82_ab_29__23_, u5_mult_82_ab_29__24_, u5_mult_82_ab_29__25_,
         u5_mult_82_ab_29__26_, u5_mult_82_ab_29__27_, u5_mult_82_ab_29__28_,
         u5_mult_82_ab_29__29_, u5_mult_82_ab_29__30_, u5_mult_82_ab_29__31_,
         u5_mult_82_ab_29__32_, u5_mult_82_ab_29__33_, u5_mult_82_ab_29__34_,
         u5_mult_82_ab_29__35_, u5_mult_82_ab_29__36_, u5_mult_82_ab_29__37_,
         u5_mult_82_ab_29__38_, u5_mult_82_ab_29__39_, u5_mult_82_ab_29__40_,
         u5_mult_82_ab_29__41_, u5_mult_82_ab_29__42_, u5_mult_82_ab_29__43_,
         u5_mult_82_ab_29__44_, u5_mult_82_ab_29__45_, u5_mult_82_ab_29__46_,
         u5_mult_82_ab_29__47_, u5_mult_82_ab_29__48_, u5_mult_82_ab_29__49_,
         u5_mult_82_ab_29__50_, u5_mult_82_ab_29__51_, u5_mult_82_ab_29__52_,
         u5_mult_82_ab_30__0_, u5_mult_82_ab_30__1_, u5_mult_82_ab_30__2_,
         u5_mult_82_ab_30__3_, u5_mult_82_ab_30__4_, u5_mult_82_ab_30__5_,
         u5_mult_82_ab_30__6_, u5_mult_82_ab_30__7_, u5_mult_82_ab_30__8_,
         u5_mult_82_ab_30__9_, u5_mult_82_ab_30__10_, u5_mult_82_ab_30__11_,
         u5_mult_82_ab_30__12_, u5_mult_82_ab_30__13_, u5_mult_82_ab_30__14_,
         u5_mult_82_ab_30__15_, u5_mult_82_ab_30__16_, u5_mult_82_ab_30__17_,
         u5_mult_82_ab_30__18_, u5_mult_82_ab_30__19_, u5_mult_82_ab_30__20_,
         u5_mult_82_ab_30__21_, u5_mult_82_ab_30__22_, u5_mult_82_ab_30__23_,
         u5_mult_82_ab_30__24_, u5_mult_82_ab_30__25_, u5_mult_82_ab_30__26_,
         u5_mult_82_ab_30__27_, u5_mult_82_ab_30__28_, u5_mult_82_ab_30__29_,
         u5_mult_82_ab_30__30_, u5_mult_82_ab_30__31_, u5_mult_82_ab_30__32_,
         u5_mult_82_ab_30__33_, u5_mult_82_ab_30__34_, u5_mult_82_ab_30__35_,
         u5_mult_82_ab_30__36_, u5_mult_82_ab_30__37_, u5_mult_82_ab_30__38_,
         u5_mult_82_ab_30__39_, u5_mult_82_ab_30__40_, u5_mult_82_ab_30__41_,
         u5_mult_82_ab_30__42_, u5_mult_82_ab_30__43_, u5_mult_82_ab_30__44_,
         u5_mult_82_ab_30__45_, u5_mult_82_ab_30__46_, u5_mult_82_ab_30__47_,
         u5_mult_82_ab_30__48_, u5_mult_82_ab_30__49_, u5_mult_82_ab_30__50_,
         u5_mult_82_ab_30__51_, u5_mult_82_ab_30__52_, u5_mult_82_ab_31__0_,
         u5_mult_82_ab_31__1_, u5_mult_82_ab_31__2_, u5_mult_82_ab_31__3_,
         u5_mult_82_ab_31__4_, u5_mult_82_ab_31__5_, u5_mult_82_ab_31__6_,
         u5_mult_82_ab_31__7_, u5_mult_82_ab_31__8_, u5_mult_82_ab_31__9_,
         u5_mult_82_ab_31__10_, u5_mult_82_ab_31__11_, u5_mult_82_ab_31__12_,
         u5_mult_82_ab_31__13_, u5_mult_82_ab_31__14_, u5_mult_82_ab_31__15_,
         u5_mult_82_ab_31__16_, u5_mult_82_ab_31__17_, u5_mult_82_ab_31__18_,
         u5_mult_82_ab_31__19_, u5_mult_82_ab_31__20_, u5_mult_82_ab_31__21_,
         u5_mult_82_ab_31__22_, u5_mult_82_ab_31__23_, u5_mult_82_ab_31__24_,
         u5_mult_82_ab_31__25_, u5_mult_82_ab_31__26_, u5_mult_82_ab_31__27_,
         u5_mult_82_ab_31__28_, u5_mult_82_ab_31__29_, u5_mult_82_ab_31__30_,
         u5_mult_82_ab_31__31_, u5_mult_82_ab_31__32_, u5_mult_82_ab_31__33_,
         u5_mult_82_ab_31__34_, u5_mult_82_ab_31__35_, u5_mult_82_ab_31__36_,
         u5_mult_82_ab_31__37_, u5_mult_82_ab_31__38_, u5_mult_82_ab_31__39_,
         u5_mult_82_ab_31__40_, u5_mult_82_ab_31__41_, u5_mult_82_ab_31__42_,
         u5_mult_82_ab_31__43_, u5_mult_82_ab_31__44_, u5_mult_82_ab_31__45_,
         u5_mult_82_ab_31__46_, u5_mult_82_ab_31__47_, u5_mult_82_ab_31__48_,
         u5_mult_82_ab_31__49_, u5_mult_82_ab_31__50_, u5_mult_82_ab_31__51_,
         u5_mult_82_ab_31__52_, u5_mult_82_ab_32__0_, u5_mult_82_ab_32__1_,
         u5_mult_82_ab_32__2_, u5_mult_82_ab_32__3_, u5_mult_82_ab_32__4_,
         u5_mult_82_ab_32__5_, u5_mult_82_ab_32__6_, u5_mult_82_ab_32__7_,
         u5_mult_82_ab_32__8_, u5_mult_82_ab_32__9_, u5_mult_82_ab_32__10_,
         u5_mult_82_ab_32__11_, u5_mult_82_ab_32__12_, u5_mult_82_ab_32__13_,
         u5_mult_82_ab_32__14_, u5_mult_82_ab_32__15_, u5_mult_82_ab_32__16_,
         u5_mult_82_ab_32__17_, u5_mult_82_ab_32__18_, u5_mult_82_ab_32__19_,
         u5_mult_82_ab_32__20_, u5_mult_82_ab_32__21_, u5_mult_82_ab_32__22_,
         u5_mult_82_ab_32__23_, u5_mult_82_ab_32__24_, u5_mult_82_ab_32__25_,
         u5_mult_82_ab_32__26_, u5_mult_82_ab_32__27_, u5_mult_82_ab_32__28_,
         u5_mult_82_ab_32__29_, u5_mult_82_ab_32__30_, u5_mult_82_ab_32__31_,
         u5_mult_82_ab_32__32_, u5_mult_82_ab_32__33_, u5_mult_82_ab_32__34_,
         u5_mult_82_ab_32__35_, u5_mult_82_ab_32__36_, u5_mult_82_ab_32__37_,
         u5_mult_82_ab_32__38_, u5_mult_82_ab_32__39_, u5_mult_82_ab_32__40_,
         u5_mult_82_ab_32__41_, u5_mult_82_ab_32__42_, u5_mult_82_ab_32__43_,
         u5_mult_82_ab_32__44_, u5_mult_82_ab_32__45_, u5_mult_82_ab_32__46_,
         u5_mult_82_ab_32__47_, u5_mult_82_ab_32__48_, u5_mult_82_ab_32__49_,
         u5_mult_82_ab_32__50_, u5_mult_82_ab_32__51_, u5_mult_82_ab_32__52_,
         u5_mult_82_ab_33__0_, u5_mult_82_ab_33__1_, u5_mult_82_ab_33__2_,
         u5_mult_82_ab_33__3_, u5_mult_82_ab_33__4_, u5_mult_82_ab_33__5_,
         u5_mult_82_ab_33__6_, u5_mult_82_ab_33__7_, u5_mult_82_ab_33__8_,
         u5_mult_82_ab_33__9_, u5_mult_82_ab_33__10_, u5_mult_82_ab_33__11_,
         u5_mult_82_ab_33__12_, u5_mult_82_ab_33__13_, u5_mult_82_ab_33__14_,
         u5_mult_82_ab_33__15_, u5_mult_82_ab_33__16_, u5_mult_82_ab_33__17_,
         u5_mult_82_ab_33__18_, u5_mult_82_ab_33__19_, u5_mult_82_ab_33__20_,
         u5_mult_82_ab_33__21_, u5_mult_82_ab_33__22_, u5_mult_82_ab_33__23_,
         u5_mult_82_ab_33__24_, u5_mult_82_ab_33__25_, u5_mult_82_ab_33__26_,
         u5_mult_82_ab_33__27_, u5_mult_82_ab_33__28_, u5_mult_82_ab_33__29_,
         u5_mult_82_ab_33__30_, u5_mult_82_ab_33__31_, u5_mult_82_ab_33__32_,
         u5_mult_82_ab_33__33_, u5_mult_82_ab_33__34_, u5_mult_82_ab_33__35_,
         u5_mult_82_ab_33__36_, u5_mult_82_ab_33__37_, u5_mult_82_ab_33__38_,
         u5_mult_82_ab_33__39_, u5_mult_82_ab_33__40_, u5_mult_82_ab_33__41_,
         u5_mult_82_ab_33__42_, u5_mult_82_ab_33__43_, u5_mult_82_ab_33__44_,
         u5_mult_82_ab_33__45_, u5_mult_82_ab_33__46_, u5_mult_82_ab_33__47_,
         u5_mult_82_ab_33__48_, u5_mult_82_ab_33__49_, u5_mult_82_ab_33__50_,
         u5_mult_82_ab_33__51_, u5_mult_82_ab_33__52_, u5_mult_82_ab_34__0_,
         u5_mult_82_ab_34__1_, u5_mult_82_ab_34__2_, u5_mult_82_ab_34__3_,
         u5_mult_82_ab_34__4_, u5_mult_82_ab_34__5_, u5_mult_82_ab_34__6_,
         u5_mult_82_ab_34__7_, u5_mult_82_ab_34__8_, u5_mult_82_ab_34__9_,
         u5_mult_82_ab_34__10_, u5_mult_82_ab_34__11_, u5_mult_82_ab_34__12_,
         u5_mult_82_ab_34__13_, u5_mult_82_ab_34__14_, u5_mult_82_ab_34__15_,
         u5_mult_82_ab_34__16_, u5_mult_82_ab_34__17_, u5_mult_82_ab_34__18_,
         u5_mult_82_ab_34__19_, u5_mult_82_ab_34__20_, u5_mult_82_ab_34__21_,
         u5_mult_82_ab_34__22_, u5_mult_82_ab_34__23_, u5_mult_82_ab_34__24_,
         u5_mult_82_ab_34__25_, u5_mult_82_ab_34__26_, u5_mult_82_ab_34__27_,
         u5_mult_82_ab_34__28_, u5_mult_82_ab_34__29_, u5_mult_82_ab_34__30_,
         u5_mult_82_ab_34__31_, u5_mult_82_ab_34__32_, u5_mult_82_ab_34__33_,
         u5_mult_82_ab_34__34_, u5_mult_82_ab_34__35_, u5_mult_82_ab_34__36_,
         u5_mult_82_ab_34__37_, u5_mult_82_ab_34__38_, u5_mult_82_ab_34__39_,
         u5_mult_82_ab_34__40_, u5_mult_82_ab_34__41_, u5_mult_82_ab_34__42_,
         u5_mult_82_ab_34__43_, u5_mult_82_ab_34__44_, u5_mult_82_ab_34__45_,
         u5_mult_82_ab_34__46_, u5_mult_82_ab_34__47_, u5_mult_82_ab_34__48_,
         u5_mult_82_ab_34__49_, u5_mult_82_ab_34__50_, u5_mult_82_ab_34__51_,
         u5_mult_82_ab_34__52_, u5_mult_82_ab_35__0_, u5_mult_82_ab_35__1_,
         u5_mult_82_ab_35__2_, u5_mult_82_ab_35__3_, u5_mult_82_ab_35__4_,
         u5_mult_82_ab_35__5_, u5_mult_82_ab_35__6_, u5_mult_82_ab_35__7_,
         u5_mult_82_ab_35__8_, u5_mult_82_ab_35__9_, u5_mult_82_ab_35__10_,
         u5_mult_82_ab_35__11_, u5_mult_82_ab_35__12_, u5_mult_82_ab_35__13_,
         u5_mult_82_ab_35__14_, u5_mult_82_ab_35__15_, u5_mult_82_ab_35__16_,
         u5_mult_82_ab_35__17_, u5_mult_82_ab_35__18_, u5_mult_82_ab_35__19_,
         u5_mult_82_ab_35__20_, u5_mult_82_ab_35__21_, u5_mult_82_ab_35__22_,
         u5_mult_82_ab_35__23_, u5_mult_82_ab_35__24_, u5_mult_82_ab_35__25_,
         u5_mult_82_ab_35__26_, u5_mult_82_ab_35__27_, u5_mult_82_ab_35__28_,
         u5_mult_82_ab_35__29_, u5_mult_82_ab_35__30_, u5_mult_82_ab_35__31_,
         u5_mult_82_ab_35__32_, u5_mult_82_ab_35__33_, u5_mult_82_ab_35__34_,
         u5_mult_82_ab_35__35_, u5_mult_82_ab_35__36_, u5_mult_82_ab_35__37_,
         u5_mult_82_ab_35__38_, u5_mult_82_ab_35__39_, u5_mult_82_ab_35__40_,
         u5_mult_82_ab_35__41_, u5_mult_82_ab_35__42_, u5_mult_82_ab_35__43_,
         u5_mult_82_ab_35__44_, u5_mult_82_ab_35__45_, u5_mult_82_ab_35__46_,
         u5_mult_82_ab_35__47_, u5_mult_82_ab_35__48_, u5_mult_82_ab_35__49_,
         u5_mult_82_ab_35__50_, u5_mult_82_ab_35__51_, u5_mult_82_ab_35__52_,
         u5_mult_82_ab_36__0_, u5_mult_82_ab_36__1_, u5_mult_82_ab_36__2_,
         u5_mult_82_ab_36__3_, u5_mult_82_ab_36__4_, u5_mult_82_ab_36__5_,
         u5_mult_82_ab_36__6_, u5_mult_82_ab_36__7_, u5_mult_82_ab_36__8_,
         u5_mult_82_ab_36__9_, u5_mult_82_ab_36__10_, u5_mult_82_ab_36__11_,
         u5_mult_82_ab_36__12_, u5_mult_82_ab_36__13_, u5_mult_82_ab_36__14_,
         u5_mult_82_ab_36__15_, u5_mult_82_ab_36__16_, u5_mult_82_ab_36__17_,
         u5_mult_82_ab_36__18_, u5_mult_82_ab_36__19_, u5_mult_82_ab_36__20_,
         u5_mult_82_ab_36__21_, u5_mult_82_ab_36__22_, u5_mult_82_ab_36__23_,
         u5_mult_82_ab_36__24_, u5_mult_82_ab_36__25_, u5_mult_82_ab_36__26_,
         u5_mult_82_ab_36__27_, u5_mult_82_ab_36__28_, u5_mult_82_ab_36__29_,
         u5_mult_82_ab_36__30_, u5_mult_82_ab_36__31_, u5_mult_82_ab_36__32_,
         u5_mult_82_ab_36__33_, u5_mult_82_ab_36__34_, u5_mult_82_ab_36__35_,
         u5_mult_82_ab_36__36_, u5_mult_82_ab_36__37_, u5_mult_82_ab_36__38_,
         u5_mult_82_ab_36__39_, u5_mult_82_ab_36__40_, u5_mult_82_ab_36__41_,
         u5_mult_82_ab_36__42_, u5_mult_82_ab_36__43_, u5_mult_82_ab_36__44_,
         u5_mult_82_ab_36__45_, u5_mult_82_ab_36__46_, u5_mult_82_ab_36__47_,
         u5_mult_82_ab_36__48_, u5_mult_82_ab_36__49_, u5_mult_82_ab_36__50_,
         u5_mult_82_ab_36__51_, u5_mult_82_ab_36__52_, u5_mult_82_ab_37__0_,
         u5_mult_82_ab_37__1_, u5_mult_82_ab_37__2_, u5_mult_82_ab_37__3_,
         u5_mult_82_ab_37__4_, u5_mult_82_ab_37__5_, u5_mult_82_ab_37__6_,
         u5_mult_82_ab_37__7_, u5_mult_82_ab_37__8_, u5_mult_82_ab_37__9_,
         u5_mult_82_ab_37__10_, u5_mult_82_ab_37__11_, u5_mult_82_ab_37__12_,
         u5_mult_82_ab_37__13_, u5_mult_82_ab_37__14_, u5_mult_82_ab_37__15_,
         u5_mult_82_ab_37__16_, u5_mult_82_ab_37__17_, u5_mult_82_ab_37__18_,
         u5_mult_82_ab_37__19_, u5_mult_82_ab_37__20_, u5_mult_82_ab_37__21_,
         u5_mult_82_ab_37__22_, u5_mult_82_ab_37__23_, u5_mult_82_ab_37__24_,
         u5_mult_82_ab_37__25_, u5_mult_82_ab_37__26_, u5_mult_82_ab_37__27_,
         u5_mult_82_ab_37__28_, u5_mult_82_ab_37__29_, u5_mult_82_ab_37__30_,
         u5_mult_82_ab_37__31_, u5_mult_82_ab_37__32_, u5_mult_82_ab_37__33_,
         u5_mult_82_ab_37__34_, u5_mult_82_ab_37__35_, u5_mult_82_ab_37__36_,
         u5_mult_82_ab_37__37_, u5_mult_82_ab_37__38_, u5_mult_82_ab_37__39_,
         u5_mult_82_ab_37__40_, u5_mult_82_ab_37__41_, u5_mult_82_ab_37__42_,
         u5_mult_82_ab_37__43_, u5_mult_82_ab_37__44_, u5_mult_82_ab_37__45_,
         u5_mult_82_ab_37__46_, u5_mult_82_ab_37__47_, u5_mult_82_ab_37__48_,
         u5_mult_82_ab_37__49_, u5_mult_82_ab_37__50_, u5_mult_82_ab_37__51_,
         u5_mult_82_ab_37__52_, u5_mult_82_ab_38__0_, u5_mult_82_ab_38__1_,
         u5_mult_82_ab_38__2_, u5_mult_82_ab_38__3_, u5_mult_82_ab_38__4_,
         u5_mult_82_ab_38__5_, u5_mult_82_ab_38__6_, u5_mult_82_ab_38__7_,
         u5_mult_82_ab_38__8_, u5_mult_82_ab_38__9_, u5_mult_82_ab_38__10_,
         u5_mult_82_ab_38__11_, u5_mult_82_ab_38__12_, u5_mult_82_ab_38__13_,
         u5_mult_82_ab_38__14_, u5_mult_82_ab_38__15_, u5_mult_82_ab_38__16_,
         u5_mult_82_ab_38__17_, u5_mult_82_ab_38__18_, u5_mult_82_ab_38__19_,
         u5_mult_82_ab_38__20_, u5_mult_82_ab_38__21_, u5_mult_82_ab_38__22_,
         u5_mult_82_ab_38__23_, u5_mult_82_ab_38__24_, u5_mult_82_ab_38__25_,
         u5_mult_82_ab_38__26_, u5_mult_82_ab_38__27_, u5_mult_82_ab_38__28_,
         u5_mult_82_ab_38__29_, u5_mult_82_ab_38__30_, u5_mult_82_ab_38__31_,
         u5_mult_82_ab_38__32_, u5_mult_82_ab_38__33_, u5_mult_82_ab_38__34_,
         u5_mult_82_ab_38__35_, u5_mult_82_ab_38__36_, u5_mult_82_ab_38__37_,
         u5_mult_82_ab_38__38_, u5_mult_82_ab_38__39_, u5_mult_82_ab_38__40_,
         u5_mult_82_ab_38__41_, u5_mult_82_ab_38__42_, u5_mult_82_ab_38__43_,
         u5_mult_82_ab_38__44_, u5_mult_82_ab_38__45_, u5_mult_82_ab_38__46_,
         u5_mult_82_ab_38__47_, u5_mult_82_ab_38__48_, u5_mult_82_ab_38__49_,
         u5_mult_82_ab_38__50_, u5_mult_82_ab_38__51_, u5_mult_82_ab_38__52_,
         u5_mult_82_ab_39__0_, u5_mult_82_ab_39__1_, u5_mult_82_ab_39__2_,
         u5_mult_82_ab_39__3_, u5_mult_82_ab_39__4_, u5_mult_82_ab_39__5_,
         u5_mult_82_ab_39__6_, u5_mult_82_ab_39__7_, u5_mult_82_ab_39__8_,
         u5_mult_82_ab_39__9_, u5_mult_82_ab_39__10_, u5_mult_82_ab_39__11_,
         u5_mult_82_ab_39__12_, u5_mult_82_ab_39__13_, u5_mult_82_ab_39__14_,
         u5_mult_82_ab_39__15_, u5_mult_82_ab_39__16_, u5_mult_82_ab_39__17_,
         u5_mult_82_ab_39__18_, u5_mult_82_ab_39__19_, u5_mult_82_ab_39__20_,
         u5_mult_82_ab_39__21_, u5_mult_82_ab_39__22_, u5_mult_82_ab_39__23_,
         u5_mult_82_ab_39__24_, u5_mult_82_ab_39__25_, u5_mult_82_ab_39__26_,
         u5_mult_82_ab_39__27_, u5_mult_82_ab_39__28_, u5_mult_82_ab_39__29_,
         u5_mult_82_ab_39__30_, u5_mult_82_ab_39__31_, u5_mult_82_ab_39__32_,
         u5_mult_82_ab_39__33_, u5_mult_82_ab_39__34_, u5_mult_82_ab_39__35_,
         u5_mult_82_ab_39__36_, u5_mult_82_ab_39__37_, u5_mult_82_ab_39__38_,
         u5_mult_82_ab_39__39_, u5_mult_82_ab_39__40_, u5_mult_82_ab_39__41_,
         u5_mult_82_ab_39__42_, u5_mult_82_ab_39__43_, u5_mult_82_ab_39__44_,
         u5_mult_82_ab_39__45_, u5_mult_82_ab_39__46_, u5_mult_82_ab_39__47_,
         u5_mult_82_ab_39__48_, u5_mult_82_ab_39__49_, u5_mult_82_ab_39__50_,
         u5_mult_82_ab_39__51_, u5_mult_82_ab_39__52_, u5_mult_82_ab_40__0_,
         u5_mult_82_ab_40__1_, u5_mult_82_ab_40__2_, u5_mult_82_ab_40__3_,
         u5_mult_82_ab_40__4_, u5_mult_82_ab_40__5_, u5_mult_82_ab_40__6_,
         u5_mult_82_ab_40__7_, u5_mult_82_ab_40__8_, u5_mult_82_ab_40__9_,
         u5_mult_82_ab_40__10_, u5_mult_82_ab_40__11_, u5_mult_82_ab_40__12_,
         u5_mult_82_ab_40__13_, u5_mult_82_ab_40__14_, u5_mult_82_ab_40__15_,
         u5_mult_82_ab_40__16_, u5_mult_82_ab_40__17_, u5_mult_82_ab_40__18_,
         u5_mult_82_ab_40__19_, u5_mult_82_ab_40__20_, u5_mult_82_ab_40__21_,
         u5_mult_82_ab_40__22_, u5_mult_82_ab_40__23_, u5_mult_82_ab_40__24_,
         u5_mult_82_ab_40__25_, u5_mult_82_ab_40__26_, u5_mult_82_ab_40__27_,
         u5_mult_82_ab_40__28_, u5_mult_82_ab_40__29_, u5_mult_82_ab_40__30_,
         u5_mult_82_ab_40__31_, u5_mult_82_ab_40__32_, u5_mult_82_ab_40__33_,
         u5_mult_82_ab_40__34_, u5_mult_82_ab_40__35_, u5_mult_82_ab_40__36_,
         u5_mult_82_ab_40__37_, u5_mult_82_ab_40__38_, u5_mult_82_ab_40__39_,
         u5_mult_82_ab_40__40_, u5_mult_82_ab_40__41_, u5_mult_82_ab_40__42_,
         u5_mult_82_ab_40__43_, u5_mult_82_ab_40__44_, u5_mult_82_ab_40__45_,
         u5_mult_82_ab_40__46_, u5_mult_82_ab_40__47_, u5_mult_82_ab_40__48_,
         u5_mult_82_ab_40__49_, u5_mult_82_ab_40__50_, u5_mult_82_ab_40__51_,
         u5_mult_82_ab_40__52_, u5_mult_82_ab_41__0_, u5_mult_82_ab_41__1_,
         u5_mult_82_ab_41__2_, u5_mult_82_ab_41__3_, u5_mult_82_ab_41__4_,
         u5_mult_82_ab_41__5_, u5_mult_82_ab_41__6_, u5_mult_82_ab_41__7_,
         u5_mult_82_ab_41__8_, u5_mult_82_ab_41__9_, u5_mult_82_ab_41__10_,
         u5_mult_82_ab_41__11_, u5_mult_82_ab_41__12_, u5_mult_82_ab_41__13_,
         u5_mult_82_ab_41__14_, u5_mult_82_ab_41__15_, u5_mult_82_ab_41__16_,
         u5_mult_82_ab_41__17_, u5_mult_82_ab_41__18_, u5_mult_82_ab_41__19_,
         u5_mult_82_ab_41__20_, u5_mult_82_ab_41__21_, u5_mult_82_ab_41__22_,
         u5_mult_82_ab_41__23_, u5_mult_82_ab_41__24_, u5_mult_82_ab_41__25_,
         u5_mult_82_ab_41__26_, u5_mult_82_ab_41__27_, u5_mult_82_ab_41__28_,
         u5_mult_82_ab_41__29_, u5_mult_82_ab_41__30_, u5_mult_82_ab_41__31_,
         u5_mult_82_ab_41__32_, u5_mult_82_ab_41__33_, u5_mult_82_ab_41__34_,
         u5_mult_82_ab_41__35_, u5_mult_82_ab_41__36_, u5_mult_82_ab_41__37_,
         u5_mult_82_ab_41__38_, u5_mult_82_ab_41__39_, u5_mult_82_ab_41__40_,
         u5_mult_82_ab_41__41_, u5_mult_82_ab_41__42_, u5_mult_82_ab_41__43_,
         u5_mult_82_ab_41__44_, u5_mult_82_ab_41__45_, u5_mult_82_ab_41__46_,
         u5_mult_82_ab_41__47_, u5_mult_82_ab_41__48_, u5_mult_82_ab_41__49_,
         u5_mult_82_ab_41__50_, u5_mult_82_ab_41__51_, u5_mult_82_ab_41__52_,
         u5_mult_82_ab_42__0_, u5_mult_82_ab_42__1_, u5_mult_82_ab_42__2_,
         u5_mult_82_ab_42__3_, u5_mult_82_ab_42__4_, u5_mult_82_ab_42__5_,
         u5_mult_82_ab_42__6_, u5_mult_82_ab_42__7_, u5_mult_82_ab_42__8_,
         u5_mult_82_ab_42__9_, u5_mult_82_ab_42__10_, u5_mult_82_ab_42__11_,
         u5_mult_82_ab_42__12_, u5_mult_82_ab_42__13_, u5_mult_82_ab_42__14_,
         u5_mult_82_ab_42__15_, u5_mult_82_ab_42__16_, u5_mult_82_ab_42__17_,
         u5_mult_82_ab_42__18_, u5_mult_82_ab_42__19_, u5_mult_82_ab_42__20_,
         u5_mult_82_ab_42__21_, u5_mult_82_ab_42__22_, u5_mult_82_ab_42__23_,
         u5_mult_82_ab_42__24_, u5_mult_82_ab_42__25_, u5_mult_82_ab_42__26_,
         u5_mult_82_ab_42__27_, u5_mult_82_ab_42__28_, u5_mult_82_ab_42__29_,
         u5_mult_82_ab_42__30_, u5_mult_82_ab_42__31_, u5_mult_82_ab_42__32_,
         u5_mult_82_ab_42__33_, u5_mult_82_ab_42__34_, u5_mult_82_ab_42__35_,
         u5_mult_82_ab_42__36_, u5_mult_82_ab_42__37_, u5_mult_82_ab_42__38_,
         u5_mult_82_ab_42__39_, u5_mult_82_ab_42__40_, u5_mult_82_ab_42__41_,
         u5_mult_82_ab_42__42_, u5_mult_82_ab_42__43_, u5_mult_82_ab_42__44_,
         u5_mult_82_ab_42__45_, u5_mult_82_ab_42__46_, u5_mult_82_ab_42__47_,
         u5_mult_82_ab_42__48_, u5_mult_82_ab_42__49_, u5_mult_82_ab_42__50_,
         u5_mult_82_ab_42__51_, u5_mult_82_ab_42__52_, u5_mult_82_ab_43__0_,
         u5_mult_82_ab_43__1_, u5_mult_82_ab_43__2_, u5_mult_82_ab_43__3_,
         u5_mult_82_ab_43__4_, u5_mult_82_ab_43__5_, u5_mult_82_ab_43__6_,
         u5_mult_82_ab_43__7_, u5_mult_82_ab_43__8_, u5_mult_82_ab_43__9_,
         u5_mult_82_ab_43__10_, u5_mult_82_ab_43__11_, u5_mult_82_ab_43__12_,
         u5_mult_82_ab_43__13_, u5_mult_82_ab_43__14_, u5_mult_82_ab_43__15_,
         u5_mult_82_ab_43__16_, u5_mult_82_ab_43__17_, u5_mult_82_ab_43__18_,
         u5_mult_82_ab_43__19_, u5_mult_82_ab_43__20_, u5_mult_82_ab_43__21_,
         u5_mult_82_ab_43__22_, u5_mult_82_ab_43__23_, u5_mult_82_ab_43__24_,
         u5_mult_82_ab_43__25_, u5_mult_82_ab_43__26_, u5_mult_82_ab_43__27_,
         u5_mult_82_ab_43__28_, u5_mult_82_ab_43__29_, u5_mult_82_ab_43__30_,
         u5_mult_82_ab_43__31_, u5_mult_82_ab_43__32_, u5_mult_82_ab_43__33_,
         u5_mult_82_ab_43__34_, u5_mult_82_ab_43__35_, u5_mult_82_ab_43__36_,
         u5_mult_82_ab_43__37_, u5_mult_82_ab_43__38_, u5_mult_82_ab_43__39_,
         u5_mult_82_ab_43__40_, u5_mult_82_ab_43__41_, u5_mult_82_ab_43__42_,
         u5_mult_82_ab_43__43_, u5_mult_82_ab_43__44_, u5_mult_82_ab_43__45_,
         u5_mult_82_ab_43__46_, u5_mult_82_ab_43__47_, u5_mult_82_ab_43__48_,
         u5_mult_82_ab_43__49_, u5_mult_82_ab_43__50_, u5_mult_82_ab_43__51_,
         u5_mult_82_ab_43__52_, u5_mult_82_ab_44__0_, u5_mult_82_ab_44__1_,
         u5_mult_82_ab_44__2_, u5_mult_82_ab_44__3_, u5_mult_82_ab_44__4_,
         u5_mult_82_ab_44__5_, u5_mult_82_ab_44__6_, u5_mult_82_ab_44__7_,
         u5_mult_82_ab_44__8_, u5_mult_82_ab_44__9_, u5_mult_82_ab_44__10_,
         u5_mult_82_ab_44__11_, u5_mult_82_ab_44__12_, u5_mult_82_ab_44__13_,
         u5_mult_82_ab_44__14_, u5_mult_82_ab_44__15_, u5_mult_82_ab_44__16_,
         u5_mult_82_ab_44__17_, u5_mult_82_ab_44__18_, u5_mult_82_ab_44__19_,
         u5_mult_82_ab_44__20_, u5_mult_82_ab_44__21_, u5_mult_82_ab_44__22_,
         u5_mult_82_ab_44__23_, u5_mult_82_ab_44__24_, u5_mult_82_ab_44__25_,
         u5_mult_82_ab_44__26_, u5_mult_82_ab_44__27_, u5_mult_82_ab_44__28_,
         u5_mult_82_ab_44__29_, u5_mult_82_ab_44__30_, u5_mult_82_ab_44__31_,
         u5_mult_82_ab_44__32_, u5_mult_82_ab_44__33_, u5_mult_82_ab_44__34_,
         u5_mult_82_ab_44__35_, u5_mult_82_ab_44__36_, u5_mult_82_ab_44__37_,
         u5_mult_82_ab_44__38_, u5_mult_82_ab_44__39_, u5_mult_82_ab_44__40_,
         u5_mult_82_ab_44__41_, u5_mult_82_ab_44__42_, u5_mult_82_ab_44__43_,
         u5_mult_82_ab_44__44_, u5_mult_82_ab_44__45_, u5_mult_82_ab_44__46_,
         u5_mult_82_ab_44__47_, u5_mult_82_ab_44__48_, u5_mult_82_ab_44__49_,
         u5_mult_82_ab_44__50_, u5_mult_82_ab_44__51_, u5_mult_82_ab_44__52_,
         u5_mult_82_ab_45__0_, u5_mult_82_ab_45__1_, u5_mult_82_ab_45__2_,
         u5_mult_82_ab_45__3_, u5_mult_82_ab_45__4_, u5_mult_82_ab_45__5_,
         u5_mult_82_ab_45__6_, u5_mult_82_ab_45__7_, u5_mult_82_ab_45__8_,
         u5_mult_82_ab_45__9_, u5_mult_82_ab_45__10_, u5_mult_82_ab_45__11_,
         u5_mult_82_ab_45__12_, u5_mult_82_ab_45__13_, u5_mult_82_ab_45__14_,
         u5_mult_82_ab_45__15_, u5_mult_82_ab_45__16_, u5_mult_82_ab_45__17_,
         u5_mult_82_ab_45__18_, u5_mult_82_ab_45__19_, u5_mult_82_ab_45__20_,
         u5_mult_82_ab_45__21_, u5_mult_82_ab_45__22_, u5_mult_82_ab_45__23_,
         u5_mult_82_ab_45__24_, u5_mult_82_ab_45__25_, u5_mult_82_ab_45__26_,
         u5_mult_82_ab_45__27_, u5_mult_82_ab_45__28_, u5_mult_82_ab_45__29_,
         u5_mult_82_ab_45__30_, u5_mult_82_ab_45__31_, u5_mult_82_ab_45__32_,
         u5_mult_82_ab_45__33_, u5_mult_82_ab_45__34_, u5_mult_82_ab_45__35_,
         u5_mult_82_ab_45__36_, u5_mult_82_ab_45__37_, u5_mult_82_ab_45__38_,
         u5_mult_82_ab_45__39_, u5_mult_82_ab_45__40_, u5_mult_82_ab_45__41_,
         u5_mult_82_ab_45__42_, u5_mult_82_ab_45__43_, u5_mult_82_ab_45__44_,
         u5_mult_82_ab_45__45_, u5_mult_82_ab_45__46_, u5_mult_82_ab_45__47_,
         u5_mult_82_ab_45__48_, u5_mult_82_ab_45__49_, u5_mult_82_ab_45__50_,
         u5_mult_82_ab_45__51_, u5_mult_82_ab_45__52_, u5_mult_82_ab_46__0_,
         u5_mult_82_ab_46__1_, u5_mult_82_ab_46__2_, u5_mult_82_ab_46__3_,
         u5_mult_82_ab_46__4_, u5_mult_82_ab_46__5_, u5_mult_82_ab_46__6_,
         u5_mult_82_ab_46__7_, u5_mult_82_ab_46__8_, u5_mult_82_ab_46__9_,
         u5_mult_82_ab_46__10_, u5_mult_82_ab_46__11_, u5_mult_82_ab_46__12_,
         u5_mult_82_ab_46__13_, u5_mult_82_ab_46__14_, u5_mult_82_ab_46__15_,
         u5_mult_82_ab_46__16_, u5_mult_82_ab_46__17_, u5_mult_82_ab_46__18_,
         u5_mult_82_ab_46__19_, u5_mult_82_ab_46__20_, u5_mult_82_ab_46__21_,
         u5_mult_82_ab_46__22_, u5_mult_82_ab_46__23_, u5_mult_82_ab_46__24_,
         u5_mult_82_ab_46__25_, u5_mult_82_ab_46__26_, u5_mult_82_ab_46__27_,
         u5_mult_82_ab_46__28_, u5_mult_82_ab_46__29_, u5_mult_82_ab_46__30_,
         u5_mult_82_ab_46__31_, u5_mult_82_ab_46__32_, u5_mult_82_ab_46__33_,
         u5_mult_82_ab_46__34_, u5_mult_82_ab_46__35_, u5_mult_82_ab_46__36_,
         u5_mult_82_ab_46__37_, u5_mult_82_ab_46__38_, u5_mult_82_ab_46__39_,
         u5_mult_82_ab_46__40_, u5_mult_82_ab_46__41_, u5_mult_82_ab_46__42_,
         u5_mult_82_ab_46__43_, u5_mult_82_ab_46__44_, u5_mult_82_ab_46__45_,
         u5_mult_82_ab_46__46_, u5_mult_82_ab_46__47_, u5_mult_82_ab_46__48_,
         u5_mult_82_ab_46__49_, u5_mult_82_ab_46__50_, u5_mult_82_ab_46__51_,
         u5_mult_82_ab_46__52_, u5_mult_82_ab_47__0_, u5_mult_82_ab_47__1_,
         u5_mult_82_ab_47__2_, u5_mult_82_ab_47__3_, u5_mult_82_ab_47__4_,
         u5_mult_82_ab_47__5_, u5_mult_82_ab_47__6_, u5_mult_82_ab_47__7_,
         u5_mult_82_ab_47__8_, u5_mult_82_ab_47__9_, u5_mult_82_ab_47__10_,
         u5_mult_82_ab_47__11_, u5_mult_82_ab_47__12_, u5_mult_82_ab_47__13_,
         u5_mult_82_ab_47__14_, u5_mult_82_ab_47__15_, u5_mult_82_ab_47__16_,
         u5_mult_82_ab_47__17_, u5_mult_82_ab_47__18_, u5_mult_82_ab_47__19_,
         u5_mult_82_ab_47__20_, u5_mult_82_ab_47__21_, u5_mult_82_ab_47__22_,
         u5_mult_82_ab_47__23_, u5_mult_82_ab_47__24_, u5_mult_82_ab_47__25_,
         u5_mult_82_ab_47__26_, u5_mult_82_ab_47__27_, u5_mult_82_ab_47__28_,
         u5_mult_82_ab_47__29_, u5_mult_82_ab_47__30_, u5_mult_82_ab_47__31_,
         u5_mult_82_ab_47__32_, u5_mult_82_ab_47__33_, u5_mult_82_ab_47__34_,
         u5_mult_82_ab_47__35_, u5_mult_82_ab_47__36_, u5_mult_82_ab_47__37_,
         u5_mult_82_ab_47__38_, u5_mult_82_ab_47__39_, u5_mult_82_ab_47__40_,
         u5_mult_82_ab_47__41_, u5_mult_82_ab_47__42_, u5_mult_82_ab_47__43_,
         u5_mult_82_ab_47__44_, u5_mult_82_ab_47__45_, u5_mult_82_ab_47__46_,
         u5_mult_82_ab_47__47_, u5_mult_82_ab_47__48_, u5_mult_82_ab_47__49_,
         u5_mult_82_ab_47__50_, u5_mult_82_ab_47__51_, u5_mult_82_ab_47__52_,
         u5_mult_82_ab_48__0_, u5_mult_82_ab_48__1_, u5_mult_82_ab_48__2_,
         u5_mult_82_ab_48__3_, u5_mult_82_ab_48__4_, u5_mult_82_ab_48__5_,
         u5_mult_82_ab_48__6_, u5_mult_82_ab_48__7_, u5_mult_82_ab_48__8_,
         u5_mult_82_ab_48__9_, u5_mult_82_ab_48__10_, u5_mult_82_ab_48__11_,
         u5_mult_82_ab_48__12_, u5_mult_82_ab_48__13_, u5_mult_82_ab_48__14_,
         u5_mult_82_ab_48__15_, u5_mult_82_ab_48__16_, u5_mult_82_ab_48__17_,
         u5_mult_82_ab_48__18_, u5_mult_82_ab_48__19_, u5_mult_82_ab_48__20_,
         u5_mult_82_ab_48__21_, u5_mult_82_ab_48__22_, u5_mult_82_ab_48__23_,
         u5_mult_82_ab_48__24_, u5_mult_82_ab_48__25_, u5_mult_82_ab_48__26_,
         u5_mult_82_ab_48__27_, u5_mult_82_ab_48__28_, u5_mult_82_ab_48__29_,
         u5_mult_82_ab_48__30_, u5_mult_82_ab_48__31_, u5_mult_82_ab_48__32_,
         u5_mult_82_ab_48__33_, u5_mult_82_ab_48__34_, u5_mult_82_ab_48__35_,
         u5_mult_82_ab_48__36_, u5_mult_82_ab_48__37_, u5_mult_82_ab_48__38_,
         u5_mult_82_ab_48__39_, u5_mult_82_ab_48__40_, u5_mult_82_ab_48__41_,
         u5_mult_82_ab_48__42_, u5_mult_82_ab_48__43_, u5_mult_82_ab_48__44_,
         u5_mult_82_ab_48__45_, u5_mult_82_ab_48__46_, u5_mult_82_ab_48__47_,
         u5_mult_82_ab_48__48_, u5_mult_82_ab_48__49_, u5_mult_82_ab_48__50_,
         u5_mult_82_ab_48__51_, u5_mult_82_ab_48__52_, u5_mult_82_ab_49__0_,
         u5_mult_82_ab_49__1_, u5_mult_82_ab_49__2_, u5_mult_82_ab_49__3_,
         u5_mult_82_ab_49__4_, u5_mult_82_ab_49__5_, u5_mult_82_ab_49__6_,
         u5_mult_82_ab_49__7_, u5_mult_82_ab_49__8_, u5_mult_82_ab_49__9_,
         u5_mult_82_ab_49__10_, u5_mult_82_ab_49__11_, u5_mult_82_ab_49__12_,
         u5_mult_82_ab_49__13_, u5_mult_82_ab_49__14_, u5_mult_82_ab_49__15_,
         u5_mult_82_ab_49__16_, u5_mult_82_ab_49__17_, u5_mult_82_ab_49__18_,
         u5_mult_82_ab_49__19_, u5_mult_82_ab_49__20_, u5_mult_82_ab_49__21_,
         u5_mult_82_ab_49__22_, u5_mult_82_ab_49__23_, u5_mult_82_ab_49__24_,
         u5_mult_82_ab_49__25_, u5_mult_82_ab_49__26_, u5_mult_82_ab_49__27_,
         u5_mult_82_ab_49__28_, u5_mult_82_ab_49__29_, u5_mult_82_ab_49__30_,
         u5_mult_82_ab_49__31_, u5_mult_82_ab_49__32_, u5_mult_82_ab_49__33_,
         u5_mult_82_ab_49__34_, u5_mult_82_ab_49__35_, u5_mult_82_ab_49__36_,
         u5_mult_82_ab_49__37_, u5_mult_82_ab_49__38_, u5_mult_82_ab_49__39_,
         u5_mult_82_ab_49__40_, u5_mult_82_ab_49__41_, u5_mult_82_ab_49__42_,
         u5_mult_82_ab_49__43_, u5_mult_82_ab_49__44_, u5_mult_82_ab_49__45_,
         u5_mult_82_ab_49__46_, u5_mult_82_ab_49__47_, u5_mult_82_ab_49__48_,
         u5_mult_82_ab_49__49_, u5_mult_82_ab_49__50_, u5_mult_82_ab_49__51_,
         u5_mult_82_ab_49__52_, u5_mult_82_ab_50__0_, u5_mult_82_ab_50__1_,
         u5_mult_82_ab_50__2_, u5_mult_82_ab_50__3_, u5_mult_82_ab_50__4_,
         u5_mult_82_ab_50__5_, u5_mult_82_ab_50__6_, u5_mult_82_ab_50__7_,
         u5_mult_82_ab_50__8_, u5_mult_82_ab_50__9_, u5_mult_82_ab_50__10_,
         u5_mult_82_ab_50__11_, u5_mult_82_ab_50__12_, u5_mult_82_ab_50__13_,
         u5_mult_82_ab_50__14_, u5_mult_82_ab_50__15_, u5_mult_82_ab_50__16_,
         u5_mult_82_ab_50__17_, u5_mult_82_ab_50__18_, u5_mult_82_ab_50__19_,
         u5_mult_82_ab_50__20_, u5_mult_82_ab_50__21_, u5_mult_82_ab_50__22_,
         u5_mult_82_ab_50__23_, u5_mult_82_ab_50__24_, u5_mult_82_ab_50__25_,
         u5_mult_82_ab_50__26_, u5_mult_82_ab_50__27_, u5_mult_82_ab_50__28_,
         u5_mult_82_ab_50__29_, u5_mult_82_ab_50__30_, u5_mult_82_ab_50__31_,
         u5_mult_82_ab_50__32_, u5_mult_82_ab_50__33_, u5_mult_82_ab_50__34_,
         u5_mult_82_ab_50__35_, u5_mult_82_ab_50__36_, u5_mult_82_ab_50__37_,
         u5_mult_82_ab_50__38_, u5_mult_82_ab_50__39_, u5_mult_82_ab_50__40_,
         u5_mult_82_ab_50__41_, u5_mult_82_ab_50__42_, u5_mult_82_ab_50__43_,
         u5_mult_82_ab_50__44_, u5_mult_82_ab_50__45_, u5_mult_82_ab_50__46_,
         u5_mult_82_ab_50__47_, u5_mult_82_ab_50__48_, u5_mult_82_ab_50__49_,
         u5_mult_82_ab_50__50_, u5_mult_82_ab_50__51_, u5_mult_82_ab_50__52_,
         u5_mult_82_ab_51__0_, u5_mult_82_ab_51__1_, u5_mult_82_ab_51__2_,
         u5_mult_82_ab_51__3_, u5_mult_82_ab_51__4_, u5_mult_82_ab_51__5_,
         u5_mult_82_ab_51__6_, u5_mult_82_ab_51__7_, u5_mult_82_ab_51__8_,
         u5_mult_82_ab_51__9_, u5_mult_82_ab_51__10_, u5_mult_82_ab_51__11_,
         u5_mult_82_ab_51__12_, u5_mult_82_ab_51__13_, u5_mult_82_ab_51__14_,
         u5_mult_82_ab_51__15_, u5_mult_82_ab_51__16_, u5_mult_82_ab_51__17_,
         u5_mult_82_ab_51__18_, u5_mult_82_ab_51__19_, u5_mult_82_ab_51__20_,
         u5_mult_82_ab_51__21_, u5_mult_82_ab_51__22_, u5_mult_82_ab_51__23_,
         u5_mult_82_ab_51__24_, u5_mult_82_ab_51__25_, u5_mult_82_ab_51__26_,
         u5_mult_82_ab_51__27_, u5_mult_82_ab_51__28_, u5_mult_82_ab_51__29_,
         u5_mult_82_ab_51__30_, u5_mult_82_ab_51__31_, u5_mult_82_ab_51__32_,
         u5_mult_82_ab_51__33_, u5_mult_82_ab_51__34_, u5_mult_82_ab_51__35_,
         u5_mult_82_ab_51__36_, u5_mult_82_ab_51__37_, u5_mult_82_ab_51__38_,
         u5_mult_82_ab_51__39_, u5_mult_82_ab_51__40_, u5_mult_82_ab_51__41_,
         u5_mult_82_ab_51__42_, u5_mult_82_ab_51__43_, u5_mult_82_ab_51__44_,
         u5_mult_82_ab_51__45_, u5_mult_82_ab_51__46_, u5_mult_82_ab_51__47_,
         u5_mult_82_ab_51__48_, u5_mult_82_ab_51__49_, u5_mult_82_ab_51__50_,
         u5_mult_82_ab_51__51_, u5_mult_82_ab_51__52_, u5_mult_82_ab_52__0_,
         u5_mult_82_ab_52__1_, u5_mult_82_ab_52__2_, u5_mult_82_ab_52__3_,
         u5_mult_82_ab_52__4_, u5_mult_82_ab_52__5_, u5_mult_82_ab_52__6_,
         u5_mult_82_ab_52__7_, u5_mult_82_ab_52__8_, u5_mult_82_ab_52__9_,
         u5_mult_82_ab_52__10_, u5_mult_82_ab_52__11_, u5_mult_82_ab_52__12_,
         u5_mult_82_ab_52__13_, u5_mult_82_ab_52__14_, u5_mult_82_ab_52__15_,
         u5_mult_82_ab_52__16_, u5_mult_82_ab_52__17_, u5_mult_82_ab_52__18_,
         u5_mult_82_ab_52__19_, u5_mult_82_ab_52__20_, u5_mult_82_ab_52__21_,
         u5_mult_82_ab_52__22_, u5_mult_82_ab_52__23_, u5_mult_82_ab_52__24_,
         u5_mult_82_ab_52__25_, u5_mult_82_ab_52__26_, u5_mult_82_ab_52__27_,
         u5_mult_82_ab_52__28_, u5_mult_82_ab_52__29_, u5_mult_82_ab_52__30_,
         u5_mult_82_ab_52__31_, u5_mult_82_ab_52__32_, u5_mult_82_ab_52__33_,
         u5_mult_82_ab_52__34_, u5_mult_82_ab_52__35_, u5_mult_82_ab_52__36_,
         u5_mult_82_ab_52__37_, u5_mult_82_ab_52__38_, u5_mult_82_ab_52__39_,
         u5_mult_82_ab_52__40_, u5_mult_82_ab_52__41_, u5_mult_82_ab_52__42_,
         u5_mult_82_ab_52__43_, u5_mult_82_ab_52__44_, u5_mult_82_ab_52__45_,
         u5_mult_82_ab_52__46_, u5_mult_82_ab_52__47_, u5_mult_82_ab_52__48_,
         u5_mult_82_ab_52__49_, u5_mult_82_ab_52__50_, u5_mult_82_ab_52__51_,
         u5_mult_82_ab_52__52_, u5_mult_82_FS_1_n305, u5_mult_82_FS_1_n304,
         u5_mult_82_FS_1_n303, u5_mult_82_FS_1_n302, u5_mult_82_FS_1_n301,
         u5_mult_82_FS_1_n300, u5_mult_82_FS_1_n299, u5_mult_82_FS_1_n298,
         u5_mult_82_FS_1_n297, u5_mult_82_FS_1_n296, u5_mult_82_FS_1_n295,
         u5_mult_82_FS_1_n294, u5_mult_82_FS_1_n293, u5_mult_82_FS_1_n292,
         u5_mult_82_FS_1_n291, u5_mult_82_FS_1_n290, u5_mult_82_FS_1_n289,
         u5_mult_82_FS_1_n288, u5_mult_82_FS_1_n287, u5_mult_82_FS_1_n286,
         u5_mult_82_FS_1_n285, u5_mult_82_FS_1_n284, u5_mult_82_FS_1_n283,
         u5_mult_82_FS_1_n282, u5_mult_82_FS_1_n281, u5_mult_82_FS_1_n280,
         u5_mult_82_FS_1_n279, u5_mult_82_FS_1_n278, u5_mult_82_FS_1_n277,
         u5_mult_82_FS_1_n276, u5_mult_82_FS_1_n275, u5_mult_82_FS_1_n274,
         u5_mult_82_FS_1_n273, u5_mult_82_FS_1_n272, u5_mult_82_FS_1_n271,
         u5_mult_82_FS_1_n270, u5_mult_82_FS_1_n269, u5_mult_82_FS_1_n268,
         u5_mult_82_FS_1_n267, u5_mult_82_FS_1_n266, u5_mult_82_FS_1_n265,
         u5_mult_82_FS_1_n264, u5_mult_82_FS_1_n263, u5_mult_82_FS_1_n262,
         u5_mult_82_FS_1_n261, u5_mult_82_FS_1_n260, u5_mult_82_FS_1_n259,
         u5_mult_82_FS_1_n258, u5_mult_82_FS_1_n257, u5_mult_82_FS_1_n256,
         u5_mult_82_FS_1_n255, u5_mult_82_FS_1_n254, u5_mult_82_FS_1_n253,
         u5_mult_82_FS_1_n252, u5_mult_82_FS_1_n251, u5_mult_82_FS_1_n250,
         u5_mult_82_FS_1_n249, u5_mult_82_FS_1_n248, u5_mult_82_FS_1_n247,
         u5_mult_82_FS_1_n246, u5_mult_82_FS_1_n245, u5_mult_82_FS_1_n244,
         u5_mult_82_FS_1_n243, u5_mult_82_FS_1_n242, u5_mult_82_FS_1_n241,
         u5_mult_82_FS_1_n240, u5_mult_82_FS_1_n239, u5_mult_82_FS_1_n238,
         u5_mult_82_FS_1_n237, u5_mult_82_FS_1_n236, u5_mult_82_FS_1_n235,
         u5_mult_82_FS_1_n234, u5_mult_82_FS_1_n233, u5_mult_82_FS_1_n232,
         u5_mult_82_FS_1_n231, u5_mult_82_FS_1_n230, u5_mult_82_FS_1_n229,
         u5_mult_82_FS_1_n228, u5_mult_82_FS_1_n227, u5_mult_82_FS_1_n226,
         u5_mult_82_FS_1_n225, u5_mult_82_FS_1_n224, u5_mult_82_FS_1_n223,
         u5_mult_82_FS_1_n222, u5_mult_82_FS_1_n221, u5_mult_82_FS_1_n220,
         u5_mult_82_FS_1_n219, u5_mult_82_FS_1_n218, u5_mult_82_FS_1_n217,
         u5_mult_82_FS_1_n216, u5_mult_82_FS_1_n215, u5_mult_82_FS_1_n214,
         u5_mult_82_FS_1_n213, u5_mult_82_FS_1_n212, u5_mult_82_FS_1_n211,
         u5_mult_82_FS_1_n210, u5_mult_82_FS_1_n209, u5_mult_82_FS_1_n208,
         u5_mult_82_FS_1_n207, u5_mult_82_FS_1_n206, u5_mult_82_FS_1_n205,
         u5_mult_82_FS_1_n204, u5_mult_82_FS_1_n203, u5_mult_82_FS_1_n202,
         u5_mult_82_FS_1_n201, u5_mult_82_FS_1_n200, u5_mult_82_FS_1_n199,
         u5_mult_82_FS_1_n198, u5_mult_82_FS_1_n197, u5_mult_82_FS_1_n196,
         u5_mult_82_FS_1_n195, u5_mult_82_FS_1_n194, u5_mult_82_FS_1_n193,
         u5_mult_82_FS_1_n192, u5_mult_82_FS_1_n191, u5_mult_82_FS_1_n190,
         u5_mult_82_FS_1_n189, u5_mult_82_FS_1_n188, u5_mult_82_FS_1_n187,
         u5_mult_82_FS_1_n186, u5_mult_82_FS_1_n185, u5_mult_82_FS_1_n184,
         u5_mult_82_FS_1_n183, u5_mult_82_FS_1_n182, u5_mult_82_FS_1_n181,
         u5_mult_82_FS_1_n180, u5_mult_82_FS_1_n179, u5_mult_82_FS_1_n178,
         u5_mult_82_FS_1_n177, u5_mult_82_FS_1_n176, u5_mult_82_FS_1_n175,
         u5_mult_82_FS_1_n174, u5_mult_82_FS_1_n173, u5_mult_82_FS_1_n172,
         u5_mult_82_FS_1_n171, u5_mult_82_FS_1_n170, u5_mult_82_FS_1_n169,
         u5_mult_82_FS_1_n168, u5_mult_82_FS_1_n167, u5_mult_82_FS_1_n166,
         u5_mult_82_FS_1_n165, u5_mult_82_FS_1_n164, u5_mult_82_FS_1_n163,
         u5_mult_82_FS_1_n162, u5_mult_82_FS_1_n161, u5_mult_82_FS_1_n160,
         u5_mult_82_FS_1_n159, u5_mult_82_FS_1_n158, u5_mult_82_FS_1_n157,
         u5_mult_82_FS_1_n156, u5_mult_82_FS_1_n155, u5_mult_82_FS_1_n154,
         u5_mult_82_FS_1_n153, u5_mult_82_FS_1_n152, u5_mult_82_FS_1_n151,
         u5_mult_82_FS_1_n150, u5_mult_82_FS_1_n149, u5_mult_82_FS_1_n148,
         u5_mult_82_FS_1_n147, u5_mult_82_FS_1_n146, u5_mult_82_FS_1_n145,
         u5_mult_82_FS_1_n144, u5_mult_82_FS_1_n143, u5_mult_82_FS_1_n142,
         u5_mult_82_FS_1_n141, u5_mult_82_FS_1_n140, u5_mult_82_FS_1_n139,
         u5_mult_82_FS_1_n138, u5_mult_82_FS_1_n137, u5_mult_82_FS_1_n136,
         u5_mult_82_FS_1_n135, u5_mult_82_FS_1_n134, u5_mult_82_FS_1_n133,
         u5_mult_82_FS_1_n132, u5_mult_82_FS_1_n131, u5_mult_82_FS_1_n130,
         u5_mult_82_FS_1_n129, u5_mult_82_FS_1_n128, u5_mult_82_FS_1_n127,
         u5_mult_82_FS_1_n126, u5_mult_82_FS_1_n125, u5_mult_82_FS_1_n124,
         u5_mult_82_FS_1_n123, u5_mult_82_FS_1_n122, u5_mult_82_FS_1_n121,
         u5_mult_82_FS_1_n120, u5_mult_82_FS_1_n119, u5_mult_82_FS_1_n118,
         u5_mult_82_FS_1_n117, u5_mult_82_FS_1_n116, u5_mult_82_FS_1_n115,
         u5_mult_82_FS_1_n114, u5_mult_82_FS_1_n113, u5_mult_82_FS_1_n112,
         u5_mult_82_FS_1_n111, u5_mult_82_FS_1_n110, u5_mult_82_FS_1_n109,
         u5_mult_82_FS_1_n108, u5_mult_82_FS_1_n107, u5_mult_82_FS_1_n106,
         u5_mult_82_FS_1_n105, u5_mult_82_FS_1_n104, u5_mult_82_FS_1_n103,
         u5_mult_82_FS_1_n102, u5_mult_82_FS_1_n101, u5_mult_82_FS_1_n100,
         u5_mult_82_FS_1_n99, u5_mult_82_FS_1_n98, u5_mult_82_FS_1_n97,
         u5_mult_82_FS_1_n96, u5_mult_82_FS_1_n95, u5_mult_82_FS_1_n94,
         u5_mult_82_FS_1_n93, u5_mult_82_FS_1_n92, u5_mult_82_FS_1_n91,
         u5_mult_82_FS_1_n90, u5_mult_82_FS_1_n89, u5_mult_82_FS_1_n88,
         u5_mult_82_FS_1_n87, u5_mult_82_FS_1_n86, u5_mult_82_FS_1_n85,
         u5_mult_82_FS_1_n84, u5_mult_82_FS_1_n83, u5_mult_82_FS_1_n82,
         u5_mult_82_FS_1_n81, u5_mult_82_FS_1_n80, u5_mult_82_FS_1_n79,
         u5_mult_82_FS_1_n78, u5_mult_82_FS_1_n77, u5_mult_82_FS_1_n76,
         u5_mult_82_FS_1_n75, u5_mult_82_FS_1_n74, u5_mult_82_FS_1_n73,
         u5_mult_82_FS_1_n72, u5_mult_82_FS_1_n71, u5_mult_82_FS_1_n70,
         u5_mult_82_FS_1_n69, u5_mult_82_FS_1_n68, u5_mult_82_FS_1_n67,
         u5_mult_82_FS_1_n66, u5_mult_82_FS_1_n65, u5_mult_82_FS_1_n64,
         u5_mult_82_FS_1_n63, u5_mult_82_FS_1_n62, u5_mult_82_FS_1_n61,
         u5_mult_82_FS_1_n60, u5_mult_82_FS_1_n59, u5_mult_82_FS_1_n58,
         u5_mult_82_FS_1_n57, u5_mult_82_FS_1_n56, u5_mult_82_FS_1_n55,
         u5_mult_82_FS_1_n54, u5_mult_82_FS_1_n53, u5_mult_82_FS_1_n52,
         u5_mult_82_FS_1_n51, u5_mult_82_FS_1_n50, u5_mult_82_FS_1_n49,
         u5_mult_82_FS_1_n48, u5_mult_82_FS_1_n47, u5_mult_82_FS_1_n46,
         u5_mult_82_FS_1_n45, u5_mult_82_FS_1_n44, u5_mult_82_FS_1_n43,
         u5_mult_82_FS_1_n42, u5_mult_82_FS_1_n41, u5_mult_82_FS_1_n40,
         u5_mult_82_FS_1_n39, u5_mult_82_FS_1_n38, u5_mult_82_FS_1_n37,
         u5_mult_82_FS_1_n36, u5_mult_82_FS_1_n35, u5_mult_82_FS_1_n34,
         u5_mult_82_FS_1_n33, u5_mult_82_FS_1_n32, u5_mult_82_FS_1_n31,
         u5_mult_82_FS_1_n30, u5_mult_82_FS_1_n29, u5_mult_82_FS_1_n28,
         u5_mult_82_FS_1_n27, u5_mult_82_FS_1_n26, u5_mult_82_FS_1_n25,
         u5_mult_82_FS_1_n24, u5_mult_82_FS_1_n23, u5_mult_82_FS_1_n22,
         u5_mult_82_FS_1_n21, u5_mult_82_FS_1_n20, u5_mult_82_FS_1_n19,
         u5_mult_82_FS_1_n18, u5_mult_82_FS_1_n17, u5_mult_82_FS_1_n16,
         u5_mult_82_FS_1_n15, u5_mult_82_FS_1_n14, u5_mult_82_FS_1_n13,
         u5_mult_82_FS_1_n12, u5_mult_82_FS_1_n11, u5_mult_82_FS_1_n10,
         u5_mult_82_FS_1_n9, u5_mult_82_FS_1_n8, u5_mult_82_FS_1_n7,
         u5_mult_82_FS_1_n6, u5_mult_82_FS_1_n5, u5_mult_82_FS_1_n4,
         u5_mult_82_FS_1_n3, u5_mult_82_FS_1_n1;
  wire   [63:52] opa_r;
  wire   [63:52] opb_r;
  wire   [1:0] rmode_r1;
  wire   [1:0] rmode_r2;
  wire   [1:0] rmode_r3;
  wire   [2:0] fpu_op_r1;
  wire   [2:0] fpu_op_r2;
  wire   [2:0] fpu_op_r3;
  wire   [55:0] fracta;
  wire   [55:0] fractb;
  wire   [10:0] exp_fasu;
  wire   [51:0] fracta_mul;
  wire   [7:2] exp_mul;
  wire   [1:0] exp_ovf;
  wire   [2:0] underflow_fmul_d;
  wire   [1:0] exp_ovf_r;
  wire   [56:0] fract_out_q;
  wire   [105:0] prod;
  wire   [4:0] div_opa_ldz_d;
  wire   [107:0] quo;
  wire   [107:0] remainder;
  wire   [4:0] div_opa_ldz_r1;
  wire   [4:0] div_opa_ldz_r2;
  wire   [6:1] exp_r;
  wire   [59:1] opa_r1;
  wire   [105:0] fract_i2f;
  wire   [105:50] fract_denorm;
  wire   [2:0] underflow_fmul_r;
  wire   [55:0] u1_fractb_s;
  wire   [55:0] u1_fracta_s;
  wire   [10:0] u1_exp_diff2;
  wire   [10:0] u1_exp_small;
  wire   [2:0] u2_underflow_d;
  wire   [105:0] u5_prod1;
  wire   [107:0] u6_remainder;
  wire   [107:0] u6_quo1;
  wire   [10:0] u4_div_exp3;
  wire   [117:107] u4_exp_f2i_1;
  wire   [10:0] u4_exp_fix_divb;
  wire   [10:0] u4_exp_fix_diva;
  wire   [10:0] u4_exp_out1_mi1;
  wire   [10:0] u4_exp_out_mi1;
  wire   [6:1] u4_fi_ldz_mi22;
  wire   [8:0] u4_shift_left;
  wire   [10:0] u4_shift_right;
  wire   [10:0] u4_div_shft4;
  wire   [10:2] u4_div_shft2;
  wire   [10:0] u4_div_scht1a;
  wire   [6:2] u4_sub_481_carry;
  wire   [10:1] u4_sub_412_carry;
  wire   [10:1] u4_add_411_carry;
  wire   [10:3] u4_add_410_carry;
  wire   [10:1] u4_sub_409_carry;
  wire   [6:2] u4_sub_491_carry;
  wire   [10:1] sub_1_root_sub_0_root_u4_add_497_carry;
  wire   [10:2] u4_add_464_carry;
  wire   [6:5] u4_sll_482_SHMAG;
  wire   [10:2] u4_add_466_carry;
  wire   [51:2] u4_add_396_carry;
  wire   [56:1] u3_sub_63_carry;
  wire   [55:2] u3_add_63_carry;
  wire   [10:2] u2_add_120_carry;
  wire   [10:2] u2_add_118_carry;
  wire   [10:2] u2_add_115_carry;
  wire   [11:1] u2_sub_115_carry;
  wire   [10:1] sub_1_root_u1_sub_133_aco_carry;

  OR2_X2 u4_C19042 ( .A1(u4_N6462), .A2(u4_exp_out_0_), .ZN(u4_N6463) );
  OR2_X2 u4_C19043 ( .A1(u4_N6461), .A2(u4_exp_out_1_), .ZN(u4_N6462) );
  OR2_X2 u4_C19044 ( .A1(u4_N6460), .A2(u4_exp_out_2_), .ZN(u4_N6461) );
  OR2_X2 u4_C19045 ( .A1(u4_N6459), .A2(u4_exp_out_3_), .ZN(u4_N6460) );
  OR2_X2 u4_C19046 ( .A1(u4_N6458), .A2(u4_exp_out_4_), .ZN(u4_N6459) );
  OR2_X2 u4_C19047 ( .A1(u4_N6457), .A2(u4_exp_out_5_), .ZN(u4_N6458) );
  OR2_X2 u4_C19048 ( .A1(u4_N6456), .A2(u4_exp_out_6_), .ZN(u4_N6457) );
  OR2_X2 u4_C19049 ( .A1(u4_N6455), .A2(u4_exp_out_7_), .ZN(u4_N6456) );
  OR2_X2 u4_C19050 ( .A1(u4_N6454), .A2(u4_exp_out_8_), .ZN(u4_N6455) );
  OR2_X2 u4_C19051 ( .A1(u4_exp_out_10_), .A2(u4_exp_out_9_), .ZN(u4_N6454) );
  OR2_X2 u4_C19471 ( .A1(u4_shift_right[10]), .A2(u4_shift_right[9]), .ZN(
        u4_N5904) );
  OR2_X2 u4_C19733 ( .A1(u4_N6915), .A2(u4_N6916), .ZN(u4_N6917) );
  AND2_X2 u4_C19735 ( .A1(u4_exp_out_10_), .A2(1'b1), .ZN(u4_N6916) );
  MUX2_X2 U3 ( .A(prod[105]), .B(fract_div_105_), .S(fpu_op_r3[0]), .Z(n203)
         );
  MUX2_X2 U4 ( .A(fract_out_q[56]), .B(n203), .S(fpu_op_r3[1]), .Z(n204) );
  AND2_X2 U5 ( .A1(fract_i2f[105]), .A2(n4400), .ZN(n205) );
  MUX2_X2 U6 ( .A(n204), .B(n205), .S(n4661), .Z(fract_denorm[105]) );
  NAND2_X2 U8 ( .A1(n2388), .A2(n2389), .ZN(u4_exp_out_0_) );
  NAND2_X2 U11 ( .A1(u4_div_exp3[0]), .A2(n2394), .ZN(n2396) );
  AOI22_X2 U14 ( .A1(u4_exp_f2i_1[107]), .A2(n2400), .B1(n2401), .B2(
        u4_exp_out1_0_), .ZN(n2388) );
  OAI211_X2 U15 ( .C1(n5873), .C2(n4355), .A(n2402), .B(n2403), .ZN(
        u4_exp_out_1_) );
  AOI221_X2 U16 ( .B1(u4_N6136), .B2(n2390), .C1(n2404), .C2(n6094), .A(n2405), 
        .ZN(n2403) );
  NOR2_X4 U17 ( .A1(n4653), .A2(n2399), .ZN(n2404) );
  AOI22_X2 U18 ( .A1(u4_exp_f2i_1[108]), .A2(n2400), .B1(n2401), .B2(
        u4_exp_out1_1_), .ZN(n2402) );
  OAI221_X2 U19 ( .B1(n2407), .B2(n2408), .C1(n5872), .C2(n4355), .A(n2409), 
        .ZN(u4_exp_out_2_) );
  AOI221_X2 U20 ( .B1(u4_exp_f2i_1[109]), .B2(n2400), .C1(u4_N6137), .C2(n2390), .A(n2405), .ZN(n2409) );
  OAI221_X2 U21 ( .B1(n2411), .B2(n2408), .C1(n5871), .C2(n4355), .A(n2412), 
        .ZN(u4_exp_out_3_) );
  AOI221_X2 U22 ( .B1(u4_exp_f2i_1[110]), .B2(n2400), .C1(u4_N6138), .C2(n2390), .A(n2405), .ZN(n2412) );
  OAI221_X2 U23 ( .B1(n2414), .B2(n2408), .C1(n5870), .C2(n4355), .A(n2415), 
        .ZN(u4_exp_out_4_) );
  AOI221_X2 U24 ( .B1(u4_exp_f2i_1[111]), .B2(n2400), .C1(u4_N6139), .C2(n2390), .A(n2405), .ZN(n2415) );
  OAI221_X2 U25 ( .B1(n2416), .B2(n2408), .C1(n5869), .C2(n4355), .A(n2417), 
        .ZN(u4_exp_out_5_) );
  AOI22_X2 U26 ( .A1(u4_N6140), .A2(n2390), .B1(u4_exp_f2i_1[112]), .B2(n2400), 
        .ZN(n2417) );
  OAI221_X2 U27 ( .B1(n2418), .B2(n2408), .C1(n5868), .C2(n4355), .A(n2419), 
        .ZN(u4_exp_out_6_) );
  AOI22_X2 U28 ( .A1(u4_N6141), .A2(n2390), .B1(u4_exp_f2i_1[113]), .B2(n2400), 
        .ZN(n2419) );
  OAI221_X2 U29 ( .B1(n2420), .B2(n2408), .C1(n5867), .C2(n4355), .A(n2421), 
        .ZN(u4_exp_out_7_) );
  AOI221_X2 U30 ( .B1(u4_exp_f2i_1[114]), .B2(n2400), .C1(u4_N6142), .C2(n2390), .A(n2405), .ZN(n2421) );
  AND3_X2 U31 ( .A1(opas_r2), .A2(n6343), .A3(n2422), .ZN(n2405) );
  OAI221_X2 U32 ( .B1(n2424), .B2(n2408), .C1(n5866), .C2(n4355), .A(n2425), 
        .ZN(u4_exp_out_8_) );
  OAI221_X2 U34 ( .B1(n2428), .B2(n2408), .C1(n5865), .C2(n4355), .A(n2429), 
        .ZN(u4_exp_out_9_) );
  OAI221_X2 U36 ( .B1(n2431), .B2(n2408), .C1(n5864), .C2(n4355), .A(n2432), 
        .ZN(u4_exp_out_10_) );
  OAI211_X2 U101 ( .C1(n2442), .C2(n2443), .A(n2444), .B(n2445), .ZN(
        u4_shift_right[9]) );
  AOI22_X2 U102 ( .A1(u4_div_shft2[9]), .A2(n2446), .B1(u4_exp_in_mi1_9_), 
        .B2(n2447), .ZN(n2445) );
  AOI22_X2 U103 ( .A1(u4_div_shft4[9]), .A2(n2448), .B1(u4_div_shft3_9_), .B2(
        n2449), .ZN(n2444) );
  OAI211_X2 U104 ( .C1(n2442), .C2(n2450), .A(n2451), .B(n2452), .ZN(
        u4_shift_right[8]) );
  AOI22_X2 U105 ( .A1(u4_div_shft2[8]), .A2(n2446), .B1(u4_exp_in_mi1_8_), 
        .B2(n2447), .ZN(n2452) );
  AOI22_X2 U106 ( .A1(u4_div_shft4[8]), .A2(n2448), .B1(u4_div_shft3_8_), .B2(
        n2449), .ZN(n2451) );
  OAI211_X2 U107 ( .C1(n2442), .C2(n2453), .A(n2454), .B(n2455), .ZN(
        u4_shift_right[7]) );
  AOI22_X2 U108 ( .A1(u4_div_shft2[7]), .A2(n2446), .B1(u4_exp_in_mi1_7_), 
        .B2(n2447), .ZN(n2455) );
  AOI22_X2 U109 ( .A1(u4_div_shft4[7]), .A2(n2448), .B1(u4_div_shft3_7_), .B2(
        n2449), .ZN(n2454) );
  OAI211_X2 U110 ( .C1(n2442), .C2(n2456), .A(n2457), .B(n2458), .ZN(
        u4_shift_right[6]) );
  AOI22_X2 U111 ( .A1(u4_div_shft2[6]), .A2(n2446), .B1(u4_exp_in_mi1_6_), 
        .B2(n2447), .ZN(n2458) );
  AOI22_X2 U112 ( .A1(u4_div_shft4[6]), .A2(n2448), .B1(u4_div_shft3_6_), .B2(
        n2449), .ZN(n2457) );
  OAI211_X2 U113 ( .C1(n2442), .C2(n2459), .A(n2460), .B(n2461), .ZN(
        u4_shift_right[5]) );
  AOI22_X2 U114 ( .A1(u4_div_shft2[5]), .A2(n2446), .B1(u4_exp_in_mi1_5_), 
        .B2(n2447), .ZN(n2461) );
  AOI22_X2 U115 ( .A1(u4_div_shft4[5]), .A2(n2448), .B1(u4_div_shft3_5_), .B2(
        n2449), .ZN(n2460) );
  OAI211_X2 U116 ( .C1(n2442), .C2(n2462), .A(n2463), .B(n2464), .ZN(
        u4_shift_right[4]) );
  AOI22_X2 U117 ( .A1(u4_div_shft2[4]), .A2(n2446), .B1(u4_exp_in_mi1_4_), 
        .B2(n2447), .ZN(n2464) );
  AOI22_X2 U118 ( .A1(u4_div_shft4[4]), .A2(n2448), .B1(u4_div_shft3_4_), .B2(
        n2449), .ZN(n2463) );
  OAI211_X2 U119 ( .C1(n2442), .C2(n2465), .A(n2466), .B(n2467), .ZN(
        u4_shift_right[3]) );
  AOI22_X2 U120 ( .A1(u4_div_shft2[3]), .A2(n2446), .B1(u4_exp_in_mi1_3_), 
        .B2(n2447), .ZN(n2467) );
  AOI22_X2 U121 ( .A1(u4_div_shft4[3]), .A2(n2448), .B1(u4_div_shft3_3_), .B2(
        n2449), .ZN(n2466) );
  OAI211_X2 U122 ( .C1(n2442), .C2(n2468), .A(n2469), .B(n2470), .ZN(
        u4_shift_right[2]) );
  AOI22_X2 U123 ( .A1(u4_div_shft2[2]), .A2(n2446), .B1(u4_exp_in_mi1_2_), 
        .B2(n2447), .ZN(n2470) );
  AOI22_X2 U124 ( .A1(u4_div_shft4[2]), .A2(n2448), .B1(u4_div_shft3_2_), .B2(
        n2449), .ZN(n2469) );
  OAI211_X2 U125 ( .C1(n2442), .C2(n2471), .A(n2472), .B(n2473), .ZN(
        u4_shift_right[1]) );
  AOI22_X2 U126 ( .A1(n4314), .A2(n2446), .B1(u4_exp_in_mi1_1_), .B2(n2447), 
        .ZN(n2473) );
  AOI22_X2 U127 ( .A1(u4_div_shft4[1]), .A2(n2448), .B1(u4_div_shft3_1_), .B2(
        n2449), .ZN(n2472) );
  OAI211_X2 U128 ( .C1(u4_N6915), .C2(n2442), .A(n2474), .B(n2475), .ZN(
        u4_shift_right[10]) );
  AOI22_X2 U129 ( .A1(u4_div_shft2[10]), .A2(n2446), .B1(u4_exp_in_mi1_10_), 
        .B2(n2447), .ZN(n2475) );
  AOI22_X2 U130 ( .A1(u4_div_shft4[10]), .A2(n2448), .B1(u4_div_shft3_10_), 
        .B2(n2449), .ZN(n2474) );
  OAI211_X2 U131 ( .C1(u4_exp_out_mi1[0]), .C2(n2442), .A(n2476), .B(n2477), 
        .ZN(u4_shift_right[0]) );
  AOI22_X2 U132 ( .A1(n4600), .A2(n2446), .B1(n4349), .B2(n2447), .ZN(n2477)
         );
  AOI22_X2 U134 ( .A1(u4_div_shft4[0]), .A2(n2448), .B1(u4_div_shft3_0_), .B2(
        n2449), .ZN(n2476) );
  NAND2_X2 U137 ( .A1(n2481), .A2(n2482), .ZN(u4_shift_left[8]) );
  AOI22_X2 U138 ( .A1(u4_f2i_shft_8_), .A2(n6342), .B1(n4353), .B2(n2483), 
        .ZN(n2482) );
  AOI22_X2 U139 ( .A1(u4_div_scht1a[8]), .A2(n2484), .B1(u4_exp_in_pl1_8_), 
        .B2(n2485), .ZN(n2481) );
  NAND2_X2 U140 ( .A1(n2486), .A2(n2487), .ZN(u4_shift_left[7]) );
  AOI22_X2 U141 ( .A1(u4_f2i_shft_7_), .A2(n6342), .B1(n4281), .B2(n2483), 
        .ZN(n2487) );
  AOI22_X2 U142 ( .A1(u4_div_scht1a[7]), .A2(n2484), .B1(u4_exp_in_pl1_7_), 
        .B2(n2485), .ZN(n2486) );
  INV_X4 U143 ( .A(n2488), .ZN(u4_shift_left[6]) );
  AOI221_X2 U144 ( .B1(u4_fi_ldz_6_), .B2(n2489), .C1(n2485), .C2(
        u4_exp_in_pl1_6_), .A(n2490), .ZN(n2488) );
  INV_X4 U145 ( .A(n2491), .ZN(n2490) );
  INV_X4 U147 ( .A(n2492), .ZN(u4_shift_left[5]) );
  AOI221_X2 U148 ( .B1(n2489), .B2(u4_fi_ldz_5_), .C1(n2485), .C2(
        u4_exp_in_pl1_5_), .A(n2493), .ZN(n2492) );
  INV_X4 U149 ( .A(n2494), .ZN(n2493) );
  OAI211_X2 U151 ( .C1(n2495), .C2(n6461), .A(n2496), .B(n2497), .ZN(
        u4_shift_left[4]) );
  AOI22_X2 U153 ( .A1(u4_div_scht1a[4]), .A2(n2484), .B1(u4_fi_ldz_4_), .B2(
        n2489), .ZN(n2496) );
  OAI211_X2 U154 ( .C1(n2495), .C2(n6462), .A(n2499), .B(n2500), .ZN(
        u4_shift_left[3]) );
  AOI22_X2 U156 ( .A1(u4_div_scht1a[3]), .A2(n2484), .B1(u4_fi_ldz_3_), .B2(
        n2489), .ZN(n2499) );
  OAI211_X2 U157 ( .C1(n2495), .C2(n6463), .A(n2501), .B(n2502), .ZN(
        u4_shift_left[2]) );
  AOI22_X2 U159 ( .A1(u4_div_scht1a[2]), .A2(n2484), .B1(u4_fi_ldz_2_), .B2(
        n2489), .ZN(n2501) );
  NAND2_X2 U160 ( .A1(n2503), .A2(n2504), .ZN(u4_shift_left[1]) );
  AOI221_X2 U161 ( .B1(u4_f2i_shft_1_), .B2(n6342), .C1(div_opa_ldz_r2[1]), 
        .C2(n2498), .A(n2505), .ZN(n2504) );
  INV_X4 U163 ( .A(n2511), .ZN(n2509) );
  OAI211_X2 U165 ( .C1(n2495), .C2(n4600), .A(n2512), .B(n2513), .ZN(
        u4_shift_left[0]) );
  AOI22_X2 U168 ( .A1(u4_div_scht1a[0]), .A2(n2484), .B1(u4_fi_ldz_2a_0_), 
        .B2(n2489), .ZN(n2512) );
  OAI211_X2 U169 ( .C1(n2508), .C2(n2511), .A(n2516), .B(n2517), .ZN(n2489) );
  INV_X4 U172 ( .A(n2485), .ZN(n2495) );
  INV_X4 U173 ( .A(n2519), .ZN(u4_fract_out_5_) );
  INV_X4 U174 ( .A(n2520), .ZN(u4_fract_out_51_) );
  INV_X4 U175 ( .A(n2521), .ZN(u4_fract_out_50_) );
  INV_X4 U176 ( .A(n2522), .ZN(u4_fract_out_47_) );
  INV_X4 U177 ( .A(n2523), .ZN(u4_fract_out_46_) );
  INV_X4 U178 ( .A(n2524), .ZN(u4_fract_out_45_) );
  INV_X4 U179 ( .A(n2525), .ZN(u4_fract_out_40_) );
  INV_X4 U180 ( .A(n2526), .ZN(u4_fract_out_3_) );
  INV_X4 U181 ( .A(n2527), .ZN(u4_fract_out_39_) );
  INV_X4 U182 ( .A(n2528), .ZN(u4_fract_out_35_) );
  INV_X4 U183 ( .A(n2529), .ZN(u4_fract_out_34_) );
  INV_X4 U184 ( .A(n2530), .ZN(u4_fract_out_33_) );
  INV_X4 U185 ( .A(n2531), .ZN(u4_fract_out_29_) );
  INV_X4 U186 ( .A(n2532), .ZN(u4_fract_out_28_) );
  INV_X4 U187 ( .A(n2533), .ZN(u4_fract_out_27_) );
  INV_X4 U188 ( .A(n2534), .ZN(u4_fract_out_23_) );
  INV_X4 U189 ( .A(n2535), .ZN(u4_fract_out_22_) );
  INV_X4 U190 ( .A(n2536), .ZN(u4_fract_out_21_) );
  INV_X4 U191 ( .A(n2537), .ZN(u4_fract_out_17_) );
  INV_X4 U192 ( .A(n2538), .ZN(u4_fract_out_16_) );
  INV_X4 U193 ( .A(n2539), .ZN(u4_fract_out_15_) );
  INV_X4 U194 ( .A(n2540), .ZN(u4_fract_out_11_) );
  INV_X4 U195 ( .A(n2541), .ZN(u4_fract_out_10_) );
  AND2_X2 U196 ( .A1(n2542), .A2(n6366), .ZN(u4_fi_ldz_6_) );
  NOR4_X2 U198 ( .A1(n2547), .A2(n2548), .A3(n2549), .A4(n2550), .ZN(n2546) );
  NOR4_X2 U199 ( .A1(n2551), .A2(n2552), .A3(n2553), .A4(n2554), .ZN(n2545) );
  NOR4_X2 U206 ( .A1(n2569), .A2(n2570), .A3(n2571), .A4(n6322), .ZN(n2568) );
  NAND4_X2 U208 ( .A1(n2574), .A2(n2575), .A3(n2576), .A4(n2577), .ZN(n2563)
         );
  NOR4_X2 U209 ( .A1(n2578), .A2(n2579), .A3(n2580), .A4(n2581), .ZN(n2577) );
  NOR4_X2 U210 ( .A1(n2582), .A2(n2583), .A3(n6333), .A4(n2584), .ZN(n2576) );
  NOR4_X2 U211 ( .A1(n2586), .A2(n2587), .A3(n2588), .A4(n2589), .ZN(n2575) );
  OAI211_X2 U215 ( .C1(n2593), .C2(n6328), .A(n2594), .B(n2595), .ZN(n2571) );
  OR3_X2 U221 ( .A1(n2604), .A2(n2605), .A3(n6332), .ZN(n2603) );
  NAND4_X2 U222 ( .A1(n2606), .A2(n2607), .A3(n2608), .A4(n2609), .ZN(n2569)
         );
  NOR4_X2 U223 ( .A1(n2610), .A2(n2611), .A3(n2612), .A4(n6330), .ZN(n2567) );
  NAND4_X2 U224 ( .A1(n2614), .A2(n2615), .A3(n2616), .A4(n2617), .ZN(n2610)
         );
  NOR4_X2 U225 ( .A1(n2618), .A2(n2619), .A3(n2620), .A4(n2621), .ZN(n2566) );
  NOR4_X2 U226 ( .A1(n2622), .A2(n2623), .A3(n2624), .A4(n2625), .ZN(n2565) );
  NOR4_X2 U228 ( .A1(n2583), .A2(n2611), .A3(n2630), .A4(n2631), .ZN(n2629) );
  AND3_X2 U231 ( .A1(fract_denorm[50]), .A2(n6403), .A3(n2637), .ZN(n2583) );
  AOI221_X2 U232 ( .B1(n2638), .B2(fract_denorm[98]), .C1(n2639), .C2(n6430), 
        .A(n2640), .ZN(n2628) );
  NAND4_X2 U241 ( .A1(n2655), .A2(n2656), .A3(n2657), .A4(n2658), .ZN(n2654)
         );
  NAND4_X2 U246 ( .A1(n2662), .A2(n6361), .A3(n6362), .A4(n4653), .ZN(n2656)
         );
  OR3_X2 U248 ( .A1(n2664), .A2(n2649), .A3(n2665), .ZN(n2653) );
  AND3_X2 U253 ( .A1(n2668), .A2(n6408), .A3(n2542), .ZN(n2586) );
  NAND4_X2 U256 ( .A1(n2672), .A2(n6323), .A3(n2673), .A4(n2674), .ZN(
        u4_fi_ldz_1_) );
  NOR4_X2 U257 ( .A1(n2675), .A2(n2676), .A3(n2677), .A4(n2678), .ZN(n2674) );
  OAI22_X2 U258 ( .A1(n6329), .A2(n2682), .B1(n2683), .B2(n2684), .ZN(n2675)
         );
  NAND2_X2 U259 ( .A1(n6423), .A2(n2685), .ZN(n2682) );
  OAI211_X2 U261 ( .C1(n6364), .C2(n2689), .A(n6361), .B(n6362), .ZN(n2686) );
  OR2_X2 U262 ( .A1(fract_denorm[101]), .A2(fract_denorm[102]), .ZN(n2689) );
  OR4_X2 U264 ( .A1(n2691), .A2(n2650), .A3(n6319), .A4(n2692), .ZN(n2665) );
  OR3_X2 U265 ( .A1(n2693), .A2(n2694), .A3(n2612), .ZN(n2692) );
  AND3_X2 U266 ( .A1(n2695), .A2(n6420), .A3(n2600), .ZN(n2612) );
  OR3_X2 U268 ( .A1(n2549), .A2(n2620), .A3(n2581), .ZN(n2693) );
  AND3_X2 U269 ( .A1(n2698), .A2(fract_denorm[52]), .A3(n2679), .ZN(n2581) );
  NAND4_X2 U273 ( .A1(n2602), .A2(n2702), .A3(n2703), .A4(n2704), .ZN(n2650)
         );
  AND3_X2 U275 ( .A1(n2705), .A2(fract_denorm[60]), .A3(n2562), .ZN(n2554) );
  AND3_X2 U277 ( .A1(n2706), .A2(n6406), .A3(n2542), .ZN(n2588) );
  NOR4_X2 U286 ( .A1(n6443), .A2(n2718), .A3(n2561), .A4(n6328), .ZN(n2717) );
  AOI221_X2 U289 ( .B1(n2647), .B2(fract_denorm[73]), .C1(n6336), .C2(
        fract_denorm[89]), .A(n2648), .ZN(n2713) );
  NAND4_X2 U290 ( .A1(n6321), .A2(n6320), .A3(n2719), .A4(n2720), .ZN(n2648)
         );
  AOI221_X2 U291 ( .B1(n2542), .B2(n6367), .C1(n2562), .C2(fract_denorm[65]), 
        .A(n2721), .ZN(n2720) );
  OAI221_X2 U292 ( .B1(n2593), .B2(n6328), .C1(n2722), .C2(n6332), .A(n2723), 
        .ZN(n2721) );
  AOI221_X2 U294 ( .B1(n6325), .B2(fract_denorm[81]), .C1(n6338), .C2(
        fract_denorm[97]), .A(n2701), .ZN(n2719) );
  NAND4_X2 U295 ( .A1(n2601), .A2(n2725), .A3(n2726), .A4(n2727), .ZN(n2701)
         );
  NOR4_X2 U297 ( .A1(n6334), .A2(n6388), .A3(n6387), .A4(fract_denorm[60]), 
        .ZN(n2557) );
  NAND4_X2 U298 ( .A1(n6325), .A2(n2728), .A3(fract_denorm[75]), .A4(n6381), 
        .ZN(n2617) );
  AND4_X2 U299 ( .A1(n2542), .A2(n2706), .A3(n6405), .A4(n2729), .ZN(n2589) );
  NAND4_X2 U300 ( .A1(n6338), .A2(n2707), .A3(fract_denorm[91]), .A4(n6354), 
        .ZN(n2726) );
  NAND4_X2 U301 ( .A1(n2639), .A2(n2708), .A3(n6426), .A4(n2730), .ZN(n2725)
         );
  NAND4_X2 U302 ( .A1(n2555), .A2(n2709), .A3(n6411), .A4(n2731), .ZN(n2601)
         );
  NAND4_X2 U303 ( .A1(n2606), .A2(n2732), .A3(n2733), .A4(n2734), .ZN(n2651)
         );
  AND4_X2 U305 ( .A1(n2562), .A2(n2735), .A3(fract_denorm[61]), .A4(n6389), 
        .ZN(n2553) );
  AND4_X2 U306 ( .A1(n6325), .A2(n2736), .A3(fract_denorm[77]), .A4(n6383), 
        .ZN(n2624) );
  AND4_X2 U307 ( .A1(n2542), .A2(n2668), .A3(n6407), .A4(n2737), .ZN(n2587) );
  NAND4_X2 U308 ( .A1(n6338), .A2(n2738), .A3(fract_denorm[93]), .A4(n6355), 
        .ZN(n2733) );
  NAND4_X2 U309 ( .A1(n2639), .A2(n2669), .A3(n6428), .A4(n2739), .ZN(n2732)
         );
  NAND4_X2 U310 ( .A1(n2555), .A2(n2670), .A3(n6414), .A4(n2740), .ZN(n2606)
         );
  NAND4_X2 U311 ( .A1(n2608), .A2(n2741), .A3(n2742), .A4(n2743), .ZN(n2688)
         );
  NOR4_X2 U313 ( .A1(n6334), .A2(n6392), .A3(fract_denorm[64]), .A4(
        fract_denorm[65]), .ZN(n2551) );
  NOR4_X2 U314 ( .A1(n2642), .A2(n6386), .A3(fract_denorm[80]), .A4(
        fract_denorm[81]), .ZN(n2622) );
  AND4_X2 U315 ( .A1(n2542), .A2(n6410), .A3(n2744), .A4(n2711), .ZN(n2584) );
  NAND4_X2 U316 ( .A1(n6338), .A2(fract_denorm[95]), .A3(n6356), .A4(n6358), 
        .ZN(n2742) );
  NAND4_X2 U317 ( .A1(n2639), .A2(n6432), .A3(n2681), .A4(n2722), .ZN(n2741)
         );
  NAND4_X2 U318 ( .A1(n2555), .A2(n6418), .A3(n2745), .A4(n2593), .ZN(n2608)
         );
  NAND4_X2 U321 ( .A1(n2614), .A2(n2746), .A3(n2747), .A4(n2748), .ZN(n2664)
         );
  NOR4_X2 U323 ( .A1(n6335), .A2(n6398), .A3(n6395), .A4(fract_denorm[70]), 
        .ZN(n2548) );
  AND4_X2 U324 ( .A1(n6336), .A2(n2749), .A3(fract_denorm[85]), .A4(n6376), 
        .ZN(n2619) );
  AND4_X2 U325 ( .A1(n2679), .A2(n2750), .A3(fract_denorm[53]), .A4(n6370), 
        .ZN(n2580) );
  NAND4_X2 U327 ( .A1(n6327), .A2(n2663), .A3(n6435), .A4(n2752), .ZN(n2746)
         );
  NAND4_X2 U328 ( .A1(n2600), .A2(n2660), .A3(n6421), .A4(n2753), .ZN(n2614)
         );
  NAND4_X2 U329 ( .A1(n2754), .A2(n2613), .A3(n2755), .A4(n2756), .ZN(n2691)
         );
  NOR4_X2 U330 ( .A1(n2621), .A2(n2550), .A3(n2582), .A4(n2757), .ZN(n2756) );
  NOR4_X2 U331 ( .A1(n6434), .A2(n2758), .A3(n2697), .A4(n2632), .ZN(n2757) );
  AND2_X2 U332 ( .A1(n2637), .A2(fract_denorm[51]), .ZN(n2582) );
  AND4_X2 U333 ( .A1(n2647), .A2(n2759), .A3(fract_denorm[67]), .A4(n6394), 
        .ZN(n2550) );
  AND4_X2 U334 ( .A1(n6336), .A2(n2760), .A3(fract_denorm[83]), .A4(n6374), 
        .ZN(n2621) );
  NAND4_X2 U336 ( .A1(n2600), .A2(n2695), .A3(n6419), .A4(n2762), .ZN(n2613)
         );
  NAND4_X2 U338 ( .A1(n2616), .A2(n2764), .A3(n2765), .A4(n2766), .ZN(n2690)
         );
  NOR4_X2 U340 ( .A1(n6335), .A2(n6399), .A3(fract_denorm[72]), .A4(
        fract_denorm[73]), .ZN(n2547) );
  AND4_X2 U341 ( .A1(n6336), .A2(fract_denorm[87]), .A3(n6377), .A4(n6379), 
        .ZN(n2618) );
  AND4_X2 U342 ( .A1(n2679), .A2(fract_denorm[55]), .A3(n6371), .A4(n6373), 
        .ZN(n2578) );
  OR3_X2 U343 ( .A1(n2767), .A2(n6351), .A3(n2684), .ZN(n2765) );
  NAND4_X2 U344 ( .A1(n6327), .A2(n6439), .A3(n2680), .A4(n2768), .ZN(n2764)
         );
  NAND4_X2 U345 ( .A1(n2600), .A2(n6425), .A3(n2769), .A4(n2685), .ZN(n2616)
         );
  AND3_X2 U350 ( .A1(n2698), .A2(n6400), .A3(n2679), .ZN(n2637) );
  AOI22_X2 U355 ( .A1(fract_denorm[105]), .A2(u4_exp_in_pl1_9_), .B1(n4654), 
        .B2(u4_exp_next_mi_9_), .ZN(n2428) );
  AOI22_X2 U356 ( .A1(fract_denorm[105]), .A2(u4_exp_in_pl1_8_), .B1(n4654), 
        .B2(u4_exp_next_mi_8_), .ZN(n2424) );
  AOI22_X2 U357 ( .A1(fract_denorm[105]), .A2(u4_exp_in_pl1_7_), .B1(n4654), 
        .B2(u4_exp_next_mi_7_), .ZN(n2420) );
  AOI22_X2 U358 ( .A1(fract_denorm[105]), .A2(u4_exp_in_pl1_6_), .B1(n4654), 
        .B2(u4_exp_next_mi_6_), .ZN(n2418) );
  AOI22_X2 U359 ( .A1(fract_denorm[105]), .A2(u4_exp_in_pl1_5_), .B1(n4654), 
        .B2(u4_exp_next_mi_5_), .ZN(n2416) );
  AOI22_X2 U360 ( .A1(fract_denorm[105]), .A2(u4_exp_in_pl1_4_), .B1(n4654), 
        .B2(u4_exp_next_mi_4_), .ZN(n2414) );
  AOI22_X2 U361 ( .A1(fract_denorm[105]), .A2(u4_exp_in_pl1_3_), .B1(n4654), 
        .B2(u4_exp_next_mi_3_), .ZN(n2411) );
  AOI22_X2 U362 ( .A1(fract_denorm[105]), .A2(u4_exp_in_pl1_2_), .B1(n4654), 
        .B2(u4_exp_next_mi_2_), .ZN(n2407) );
  OAI22_X2 U363 ( .A1(n4654), .A2(n6464), .B1(fract_denorm[105]), .B2(n6097), 
        .ZN(u4_exp_out1_1_) );
  AOI22_X2 U364 ( .A1(n4652), .A2(u4_exp_in_pl1_10_), .B1(n4654), .B2(
        u4_exp_next_mi_10_), .ZN(n2431) );
  OAI22_X2 U365 ( .A1(n4654), .A2(n4600), .B1(fract_denorm[105]), .B2(n6098), 
        .ZN(u4_exp_out1_0_) );
  INV_X4 U366 ( .A(u4_exp_out_10_), .ZN(u4_N6915) );
  AOI22_X2 U368 ( .A1(n2773), .A2(n2774), .B1(n2775), .B2(n2776), .ZN(n2772)
         );
  NOR4_X2 U369 ( .A1(n2777), .A2(n6034), .A3(n6036), .A4(n6035), .ZN(n2776) );
  AND4_X2 U371 ( .A1(n2779), .A2(u2_N27), .A3(u2_N25), .A4(u2_N26), .ZN(n2775)
         );
  AND3_X2 U372 ( .A1(u2_N23), .A2(u2_N22), .A3(u2_N24), .ZN(n2779) );
  NOR4_X2 U373 ( .A1(n2780), .A2(n6024), .A3(u2_N16), .A4(n4597), .ZN(n2774)
         );
  NOR4_X2 U375 ( .A1(n2781), .A2(n6026), .A3(n6030), .A4(n6028), .ZN(n2773) );
  OAI222_X2 U377 ( .A1(u6_N52), .A2(n4268), .B1(n2782), .B2(n6274), .C1(n4602), 
        .C2(n4267), .ZN(u2_underflow_d[1]) );
  AOI22_X2 U378 ( .A1(n4603), .A2(n4267), .B1(n6303), .B2(n4268), .ZN(n2783)
         );
  AND3_X2 U379 ( .A1(n6275), .A2(n2784), .A3(u2_N111), .ZN(u2_underflow_d[0])
         );
  AOI22_X2 U380 ( .A1(n4597), .A2(u2_N27), .B1(n4598), .B2(u2_N15), .ZN(n2795)
         );
  AOI22_X2 U381 ( .A1(n4597), .A2(u2_N26), .B1(n4598), .B2(u2_N14), .ZN(n2796)
         );
  AOI22_X2 U382 ( .A1(n4597), .A2(u2_N25), .B1(n4598), .B2(u2_N13), .ZN(n2797)
         );
  AOI22_X2 U383 ( .A1(n4597), .A2(u2_N24), .B1(n4598), .B2(u2_N12), .ZN(n2798)
         );
  AOI22_X2 U384 ( .A1(n4597), .A2(u2_N23), .B1(n4598), .B2(u2_N11), .ZN(n2799)
         );
  OAI22_X2 U385 ( .A1(n4599), .A2(n6033), .B1(n4597), .B2(n6024), .ZN(
        u2_exp_tmp1_4_) );
  OAI22_X2 U386 ( .A1(n4599), .A2(n6034), .B1(n4597), .B2(n6026), .ZN(
        u2_exp_tmp1_3_) );
  OAI22_X2 U387 ( .A1(n4599), .A2(n6035), .B1(n4597), .B2(n6028), .ZN(
        u2_exp_tmp1_2_) );
  OAI22_X2 U388 ( .A1(n4599), .A2(n6036), .B1(n4597), .B2(n6030), .ZN(
        u2_exp_tmp1_1_) );
  AOI22_X2 U390 ( .A1(n4597), .A2(u2_N18), .B1(n4599), .B2(u2_N6), .ZN(n2800)
         );
  OR3_X2 U392 ( .A1(n2803), .A2(n4599), .A3(n4363), .ZN(n2802) );
  NAND2_X2 U393 ( .A1(n4599), .A2(n4363), .ZN(n2801) );
  AOI22_X2 U394 ( .A1(u2_N17), .A2(n4599), .B1(u2_N29), .B2(n4597), .ZN(n2784)
         );
  OAI211_X2 U395 ( .C1(n2804), .C2(n2805), .A(n2806), .B(n2807), .ZN(u2_N86)
         );
  AOI22_X2 U396 ( .A1(u2_exp_tmp3_10_), .A2(n2808), .B1(u2_exp_tmp4_10_), .B2(
        n2809), .ZN(n2807) );
  AOI22_X2 U397 ( .A1(u2_N64), .A2(n2810), .B1(u2_N75), .B2(n2811), .ZN(n2806)
         );
  OAI211_X2 U398 ( .C1(n2785), .C2(n2805), .A(n2812), .B(n2813), .ZN(u2_N85)
         );
  AOI22_X2 U399 ( .A1(u2_exp_tmp3_9_), .A2(n2808), .B1(n2795), .B2(n2809), 
        .ZN(n2813) );
  AOI22_X2 U400 ( .A1(u2_N63), .A2(n2810), .B1(u2_N74), .B2(n2811), .ZN(n2812)
         );
  AOI22_X2 U401 ( .A1(u2_N39), .A2(n4599), .B1(u2_N51), .B2(n4597), .ZN(n2785)
         );
  OAI211_X2 U402 ( .C1(n2786), .C2(n2805), .A(n2814), .B(n2815), .ZN(u2_N84)
         );
  AOI22_X2 U403 ( .A1(u2_exp_tmp3_8_), .A2(n2808), .B1(n2796), .B2(n2809), 
        .ZN(n2815) );
  AOI22_X2 U404 ( .A1(u2_N62), .A2(n2810), .B1(u2_N73), .B2(n2811), .ZN(n2814)
         );
  AOI22_X2 U405 ( .A1(u2_N38), .A2(n4599), .B1(u2_N50), .B2(n4597), .ZN(n2786)
         );
  OAI211_X2 U406 ( .C1(n2787), .C2(n2805), .A(n2816), .B(n2817), .ZN(u2_N83)
         );
  AOI22_X2 U407 ( .A1(u2_exp_tmp3_7_), .A2(n2808), .B1(n2797), .B2(n2809), 
        .ZN(n2817) );
  AOI22_X2 U408 ( .A1(u2_N61), .A2(n2810), .B1(u2_N72), .B2(n2811), .ZN(n2816)
         );
  AOI22_X2 U409 ( .A1(u2_N37), .A2(n4599), .B1(u2_N49), .B2(n4597), .ZN(n2787)
         );
  OAI211_X2 U410 ( .C1(n2788), .C2(n2805), .A(n2818), .B(n2819), .ZN(u2_N82)
         );
  AOI22_X2 U411 ( .A1(u2_exp_tmp3_6_), .A2(n2808), .B1(n2798), .B2(n2809), 
        .ZN(n2819) );
  AOI22_X2 U412 ( .A1(u2_N60), .A2(n2810), .B1(u2_N71), .B2(n2811), .ZN(n2818)
         );
  AOI22_X2 U413 ( .A1(u2_N36), .A2(n4599), .B1(u2_N48), .B2(n4597), .ZN(n2788)
         );
  OAI211_X2 U414 ( .C1(n2789), .C2(n2805), .A(n2820), .B(n2821), .ZN(u2_N81)
         );
  AOI22_X2 U415 ( .A1(u2_exp_tmp3_5_), .A2(n2808), .B1(n2799), .B2(n2809), 
        .ZN(n2821) );
  AOI22_X2 U416 ( .A1(u2_N59), .A2(n2810), .B1(u2_N70), .B2(n2811), .ZN(n2820)
         );
  AOI22_X2 U417 ( .A1(u2_N35), .A2(n4599), .B1(u2_N47), .B2(n4597), .ZN(n2789)
         );
  OAI211_X2 U418 ( .C1(n2790), .C2(n2805), .A(n2822), .B(n2823), .ZN(u2_N80)
         );
  AOI22_X2 U419 ( .A1(u2_exp_tmp3_4_), .A2(n2808), .B1(u2_exp_tmp4_4_), .B2(
        n2809), .ZN(n2823) );
  AOI22_X2 U420 ( .A1(u2_N58), .A2(n2810), .B1(u2_N69), .B2(n2811), .ZN(n2822)
         );
  AOI22_X2 U421 ( .A1(u2_N34), .A2(n4599), .B1(u2_N46), .B2(n4597), .ZN(n2790)
         );
  OAI211_X2 U422 ( .C1(n2791), .C2(n2805), .A(n2824), .B(n2825), .ZN(u2_N79)
         );
  AOI22_X2 U423 ( .A1(u2_exp_tmp3_3_), .A2(n2808), .B1(u2_exp_tmp4_3_), .B2(
        n2809), .ZN(n2825) );
  AOI22_X2 U424 ( .A1(u2_N57), .A2(n2810), .B1(u2_N68), .B2(n2811), .ZN(n2824)
         );
  AOI22_X2 U425 ( .A1(u2_N33), .A2(n4599), .B1(u2_N45), .B2(n4597), .ZN(n2791)
         );
  OAI211_X2 U426 ( .C1(n2792), .C2(n2805), .A(n2826), .B(n2827), .ZN(u2_N78)
         );
  AOI22_X2 U427 ( .A1(u2_exp_tmp3_2_), .A2(n2808), .B1(u2_exp_tmp4_2_), .B2(
        n2809), .ZN(n2827) );
  AOI22_X2 U428 ( .A1(u2_N56), .A2(n2810), .B1(u2_N67), .B2(n2811), .ZN(n2826)
         );
  AOI22_X2 U429 ( .A1(u2_N32), .A2(n4599), .B1(u2_N44), .B2(n4597), .ZN(n2792)
         );
  OAI211_X2 U430 ( .C1(n2793), .C2(n2805), .A(n2828), .B(n2829), .ZN(u2_N77)
         );
  AOI22_X2 U431 ( .A1(u2_exp_tmp3_1_), .A2(n2808), .B1(u2_exp_tmp4_1_), .B2(
        n2809), .ZN(n2829) );
  AOI22_X2 U432 ( .A1(u2_N55), .A2(n2810), .B1(u2_N66), .B2(n2811), .ZN(n2828)
         );
  AOI22_X2 U433 ( .A1(u2_N31), .A2(n4599), .B1(u2_N43), .B2(n4597), .ZN(n2793)
         );
  OAI211_X2 U434 ( .C1(n2794), .C2(n2805), .A(n2830), .B(n2831), .ZN(u2_N76)
         );
  AOI22_X2 U435 ( .A1(u2_exp_tmp3_0_), .A2(n2808), .B1(n2800), .B2(n2809), 
        .ZN(n2831) );
  AOI22_X2 U438 ( .A1(u2_N54), .A2(n2810), .B1(u2_lt_135_A_0_), .B2(n2811), 
        .ZN(n2830) );
  NAND2_X2 U442 ( .A1(n2803), .A2(n2832), .ZN(u2_exp_ovf_d_1_) );
  AOI22_X2 U445 ( .A1(u2_N40), .A2(n4599), .B1(u2_N52), .B2(n4597), .ZN(n2804)
         );
  AOI22_X2 U446 ( .A1(u2_N41), .A2(n4599), .B1(u2_N53), .B2(n4597), .ZN(n2803)
         );
  AOI22_X2 U447 ( .A1(n2800), .A2(n4599), .B1(n2800), .B2(n4597), .ZN(n2794)
         );
  AND2_X2 U448 ( .A1(opb_r[63]), .A2(opa_r[63]), .ZN(u2_N121) );
  NAND2_X2 U450 ( .A1(u2_N113), .A2(n4597), .ZN(n2834) );
  NAND2_X2 U451 ( .A1(n6303), .A2(n4458), .ZN(n2833) );
  OAI22_X2 U453 ( .A1(n4636), .A2(n4533), .B1(n2835), .B2(n4643), .ZN(
        u1_sign_d) );
  XOR2_X2 U454 ( .A(opb_r[63]), .B(n4481), .Z(n2835) );
  OAI22_X2 U455 ( .A1(n4636), .A2(n2836), .B1(n2837), .B2(n4643), .ZN(
        u1_fractb_s[9]) );
  OAI22_X2 U456 ( .A1(n4636), .A2(n2838), .B1(n2839), .B2(n4643), .ZN(
        u1_fractb_s[8]) );
  OAI22_X2 U457 ( .A1(n4636), .A2(n2840), .B1(n2841), .B2(n4643), .ZN(
        u1_fractb_s[7]) );
  OAI22_X2 U458 ( .A1(n4636), .A2(n2842), .B1(n2843), .B2(n4643), .ZN(
        u1_fractb_s[6]) );
  OAI22_X2 U459 ( .A1(n4636), .A2(n2844), .B1(n2845), .B2(n4643), .ZN(
        u1_fractb_s[5]) );
  OAI22_X2 U460 ( .A1(n4636), .A2(n2846), .B1(n2847), .B2(n4643), .ZN(
        u1_fractb_s[55]) );
  OAI22_X2 U461 ( .A1(n4636), .A2(n2848), .B1(n2849), .B2(n4643), .ZN(
        u1_fractb_s[54]) );
  OAI22_X2 U462 ( .A1(n4636), .A2(n2850), .B1(n2851), .B2(n4643), .ZN(
        u1_fractb_s[53]) );
  OAI22_X2 U463 ( .A1(n4636), .A2(n2852), .B1(n2853), .B2(n4643), .ZN(
        u1_fractb_s[52]) );
  OAI22_X2 U464 ( .A1(n4636), .A2(n2854), .B1(n2855), .B2(n4643), .ZN(
        u1_fractb_s[51]) );
  OAI22_X2 U465 ( .A1(n4637), .A2(n2856), .B1(n2857), .B2(n4643), .ZN(
        u1_fractb_s[50]) );
  OAI22_X2 U466 ( .A1(n4637), .A2(n2858), .B1(n2859), .B2(n4643), .ZN(
        u1_fractb_s[4]) );
  OAI22_X2 U467 ( .A1(n4637), .A2(n2860), .B1(n2861), .B2(n4643), .ZN(
        u1_fractb_s[49]) );
  OAI22_X2 U468 ( .A1(n4637), .A2(n2862), .B1(n2863), .B2(n4643), .ZN(
        u1_fractb_s[48]) );
  OAI22_X2 U469 ( .A1(n4637), .A2(n2864), .B1(n2865), .B2(n4643), .ZN(
        u1_fractb_s[47]) );
  OAI22_X2 U470 ( .A1(n4637), .A2(n2866), .B1(n2867), .B2(n4643), .ZN(
        u1_fractb_s[46]) );
  OAI22_X2 U471 ( .A1(n4637), .A2(n2868), .B1(n2869), .B2(n4643), .ZN(
        u1_fractb_s[45]) );
  OAI22_X2 U472 ( .A1(n4637), .A2(n2870), .B1(n2871), .B2(n4643), .ZN(
        u1_fractb_s[44]) );
  OAI22_X2 U473 ( .A1(n4637), .A2(n2872), .B1(n2873), .B2(n4643), .ZN(
        u1_fractb_s[43]) );
  OAI22_X2 U474 ( .A1(n4637), .A2(n2874), .B1(n2875), .B2(n4643), .ZN(
        u1_fractb_s[42]) );
  OAI22_X2 U475 ( .A1(n4637), .A2(n2876), .B1(n2877), .B2(n4643), .ZN(
        u1_fractb_s[41]) );
  OAI22_X2 U476 ( .A1(n4637), .A2(n2878), .B1(n2879), .B2(n4643), .ZN(
        u1_fractb_s[40]) );
  OAI22_X2 U477 ( .A1(n4636), .A2(n2880), .B1(n2881), .B2(n4643), .ZN(
        u1_fractb_s[3]) );
  OAI22_X2 U478 ( .A1(n4639), .A2(n2882), .B1(n2883), .B2(n4644), .ZN(
        u1_fractb_s[39]) );
  OAI22_X2 U479 ( .A1(n4639), .A2(n2884), .B1(n2885), .B2(n4644), .ZN(
        u1_fractb_s[38]) );
  OAI22_X2 U480 ( .A1(n4639), .A2(n2886), .B1(n2887), .B2(n4644), .ZN(
        u1_fractb_s[37]) );
  OAI22_X2 U481 ( .A1(n4639), .A2(n2888), .B1(n2889), .B2(n4644), .ZN(
        u1_fractb_s[36]) );
  OAI22_X2 U482 ( .A1(n4639), .A2(n2890), .B1(n2891), .B2(n4644), .ZN(
        u1_fractb_s[35]) );
  OAI22_X2 U483 ( .A1(n4639), .A2(n2892), .B1(n2893), .B2(n4644), .ZN(
        u1_fractb_s[34]) );
  OAI22_X2 U484 ( .A1(n4639), .A2(n2894), .B1(n2895), .B2(n4644), .ZN(
        u1_fractb_s[33]) );
  OAI22_X2 U485 ( .A1(n4639), .A2(n2896), .B1(n2897), .B2(n4644), .ZN(
        u1_fractb_s[32]) );
  OAI22_X2 U486 ( .A1(n4639), .A2(n2898), .B1(n2899), .B2(n4644), .ZN(
        u1_fractb_s[31]) );
  OAI22_X2 U487 ( .A1(n4638), .A2(n2900), .B1(n2901), .B2(n4644), .ZN(
        u1_fractb_s[30]) );
  OAI22_X2 U488 ( .A1(n4638), .A2(n2902), .B1(n4651), .B2(n2903), .ZN(
        u1_fractb_s[2]) );
  OAI22_X2 U489 ( .A1(n4638), .A2(n2904), .B1(n2905), .B2(n4644), .ZN(
        u1_fractb_s[29]) );
  OAI22_X2 U490 ( .A1(n4638), .A2(n2906), .B1(n2907), .B2(n4644), .ZN(
        u1_fractb_s[28]) );
  OAI22_X2 U491 ( .A1(n4638), .A2(n2908), .B1(n2909), .B2(n4644), .ZN(
        u1_fractb_s[27]) );
  OAI22_X2 U492 ( .A1(n4638), .A2(n2910), .B1(n2911), .B2(n4644), .ZN(
        u1_fractb_s[26]) );
  OAI22_X2 U493 ( .A1(n4638), .A2(n2912), .B1(n2913), .B2(n4644), .ZN(
        u1_fractb_s[25]) );
  OAI22_X2 U494 ( .A1(n4638), .A2(n2914), .B1(n2915), .B2(n4644), .ZN(
        u1_fractb_s[24]) );
  OAI22_X2 U495 ( .A1(n4638), .A2(n2916), .B1(n2917), .B2(n4644), .ZN(
        u1_fractb_s[23]) );
  OAI22_X2 U496 ( .A1(n4638), .A2(n2918), .B1(n2919), .B2(n4644), .ZN(
        u1_fractb_s[22]) );
  OAI22_X2 U497 ( .A1(n4638), .A2(n2920), .B1(n2921), .B2(n4644), .ZN(
        u1_fractb_s[21]) );
  OAI22_X2 U498 ( .A1(n4639), .A2(n2922), .B1(n2923), .B2(n4644), .ZN(
        u1_fractb_s[20]) );
  OAI22_X2 U499 ( .A1(n4639), .A2(n2924), .B1(n4651), .B2(n2925), .ZN(
        u1_fractb_s[1]) );
  OAI22_X2 U500 ( .A1(n4639), .A2(n2926), .B1(n2927), .B2(n4645), .ZN(
        u1_fractb_s[19]) );
  OAI22_X2 U501 ( .A1(n4639), .A2(n2928), .B1(n2929), .B2(n4645), .ZN(
        u1_fractb_s[18]) );
  OAI22_X2 U502 ( .A1(n4639), .A2(n2930), .B1(n2931), .B2(n4645), .ZN(
        u1_fractb_s[17]) );
  OAI22_X2 U503 ( .A1(n4639), .A2(n2932), .B1(n2933), .B2(n4645), .ZN(
        u1_fractb_s[16]) );
  OAI22_X2 U504 ( .A1(n4639), .A2(n2934), .B1(n2935), .B2(n4645), .ZN(
        u1_fractb_s[15]) );
  OAI22_X2 U505 ( .A1(n4639), .A2(n2936), .B1(n2937), .B2(n4645), .ZN(
        u1_fractb_s[14]) );
  OAI22_X2 U506 ( .A1(n4639), .A2(n2938), .B1(n2939), .B2(n4645), .ZN(
        u1_fractb_s[13]) );
  OAI22_X2 U507 ( .A1(n4639), .A2(n2940), .B1(n2941), .B2(n4645), .ZN(
        u1_fractb_s[12]) );
  OAI22_X2 U508 ( .A1(n4639), .A2(n2942), .B1(n2943), .B2(n4645), .ZN(
        u1_fractb_s[11]) );
  OAI22_X2 U509 ( .A1(n4640), .A2(n2944), .B1(n2945), .B2(n4645), .ZN(
        u1_fractb_s[10]) );
  OAI22_X2 U510 ( .A1(n4640), .A2(n2946), .B1(n4651), .B2(n2947), .ZN(
        u1_fractb_s[0]) );
  OAI22_X2 U511 ( .A1(n2836), .A2(n4645), .B1(n4640), .B2(n2837), .ZN(
        u1_fracta_s[9]) );
  AOI22_X2 U512 ( .A1(n4607), .A2(u1_adj_op_out_sft_9_), .B1(n4623), .B2(u6_N6), .ZN(n2836) );
  OAI22_X2 U513 ( .A1(n2838), .A2(n4645), .B1(n4640), .B2(n2839), .ZN(
        u1_fracta_s[8]) );
  AOI22_X2 U514 ( .A1(n4606), .A2(u1_adj_op_out_sft_8_), .B1(n4621), .B2(u6_N5), .ZN(n2838) );
  OAI22_X2 U515 ( .A1(n2840), .A2(n4645), .B1(n4640), .B2(n2841), .ZN(
        u1_fracta_s[7]) );
  AOI22_X2 U516 ( .A1(n4628), .A2(u1_adj_op_out_sft_7_), .B1(n4621), .B2(u6_N4), .ZN(n2840) );
  OAI22_X2 U517 ( .A1(n2842), .A2(n4645), .B1(n4640), .B2(n2843), .ZN(
        u1_fracta_s[6]) );
  AOI22_X2 U518 ( .A1(n4615), .A2(u1_adj_op_out_sft_6_), .B1(n4621), .B2(u6_N3), .ZN(n2842) );
  OAI22_X2 U519 ( .A1(n2844), .A2(n4645), .B1(n4640), .B2(n2845), .ZN(
        u1_fracta_s[5]) );
  AOI22_X2 U520 ( .A1(n4628), .A2(u1_adj_op_out_sft_5_), .B1(n4621), .B2(u6_N2), .ZN(n2844) );
  OAI22_X2 U521 ( .A1(n2846), .A2(n4645), .B1(n4640), .B2(n2847), .ZN(
        u1_fracta_s[55]) );
  AOI22_X2 U522 ( .A1(n4606), .A2(u1_adj_op_out_sft_55_), .B1(n4621), .B2(
        u6_N52), .ZN(n2846) );
  OAI22_X2 U523 ( .A1(n2848), .A2(n4645), .B1(n4640), .B2(n2849), .ZN(
        u1_fracta_s[54]) );
  AOI22_X2 U524 ( .A1(n4606), .A2(u1_adj_op_out_sft_54_), .B1(n4621), .B2(
        u6_N51), .ZN(n2848) );
  OAI22_X2 U525 ( .A1(n2850), .A2(n4645), .B1(n4640), .B2(n2851), .ZN(
        u1_fracta_s[53]) );
  AOI22_X2 U526 ( .A1(n4606), .A2(u1_adj_op_out_sft_53_), .B1(n4621), .B2(
        u6_N50), .ZN(n2850) );
  OAI22_X2 U527 ( .A1(n2852), .A2(n4646), .B1(n4640), .B2(n2853), .ZN(
        u1_fracta_s[52]) );
  AOI22_X2 U528 ( .A1(n4606), .A2(u1_adj_op_out_sft_52_), .B1(n4621), .B2(
        u6_N49), .ZN(n2852) );
  OAI22_X2 U529 ( .A1(n2854), .A2(n4646), .B1(n4641), .B2(n2855), .ZN(
        u1_fracta_s[51]) );
  AOI22_X2 U530 ( .A1(n4606), .A2(u1_adj_op_out_sft_51_), .B1(n4621), .B2(
        u6_N48), .ZN(n2854) );
  OAI22_X2 U531 ( .A1(n2856), .A2(n4646), .B1(n4641), .B2(n2857), .ZN(
        u1_fracta_s[50]) );
  AOI22_X2 U532 ( .A1(n4606), .A2(u1_adj_op_out_sft_50_), .B1(n4621), .B2(
        u6_N47), .ZN(n2856) );
  OAI22_X2 U533 ( .A1(n2858), .A2(n4646), .B1(n4638), .B2(n2859), .ZN(
        u1_fracta_s[4]) );
  AOI22_X2 U534 ( .A1(n4628), .A2(u1_adj_op_out_sft_4_), .B1(n4621), .B2(u6_N1), .ZN(n2858) );
  OAI22_X2 U535 ( .A1(n2860), .A2(n4646), .B1(n4640), .B2(n2861), .ZN(
        u1_fracta_s[49]) );
  AOI22_X2 U536 ( .A1(n4615), .A2(u1_adj_op_out_sft_49_), .B1(n4621), .B2(
        u6_N46), .ZN(n2860) );
  OAI22_X2 U537 ( .A1(n2862), .A2(n4646), .B1(n4641), .B2(n2863), .ZN(
        u1_fracta_s[48]) );
  AOI22_X2 U538 ( .A1(n4615), .A2(u1_adj_op_out_sft_48_), .B1(n4621), .B2(
        u6_N45), .ZN(n2862) );
  OAI22_X2 U539 ( .A1(n2864), .A2(n4646), .B1(n4640), .B2(n2865), .ZN(
        u1_fracta_s[47]) );
  AOI22_X2 U540 ( .A1(n4615), .A2(u1_adj_op_out_sft_47_), .B1(n4621), .B2(
        u6_N44), .ZN(n2864) );
  OAI22_X2 U541 ( .A1(n2866), .A2(n4646), .B1(n4640), .B2(n2867), .ZN(
        u1_fracta_s[46]) );
  AOI22_X2 U542 ( .A1(n4615), .A2(u1_adj_op_out_sft_46_), .B1(n4621), .B2(
        u6_N43), .ZN(n2866) );
  OAI22_X2 U543 ( .A1(n2868), .A2(n4646), .B1(n4641), .B2(n2869), .ZN(
        u1_fracta_s[45]) );
  AOI22_X2 U544 ( .A1(n4615), .A2(u1_adj_op_out_sft_45_), .B1(n4621), .B2(
        u6_N42), .ZN(n2868) );
  OAI22_X2 U545 ( .A1(n2870), .A2(n4646), .B1(n4641), .B2(n2871), .ZN(
        u1_fracta_s[44]) );
  AOI22_X2 U546 ( .A1(n4615), .A2(u1_adj_op_out_sft_44_), .B1(n4621), .B2(
        u6_N41), .ZN(n2870) );
  OAI22_X2 U547 ( .A1(n2872), .A2(n4646), .B1(n4640), .B2(n2873), .ZN(
        u1_fracta_s[43]) );
  AOI22_X2 U548 ( .A1(n4615), .A2(u1_adj_op_out_sft_43_), .B1(n4621), .B2(
        u6_N40), .ZN(n2872) );
  OAI22_X2 U549 ( .A1(n2874), .A2(n4646), .B1(n4640), .B2(n2875), .ZN(
        u1_fracta_s[42]) );
  AOI22_X2 U550 ( .A1(n4615), .A2(u1_adj_op_out_sft_42_), .B1(n4621), .B2(
        u6_N39), .ZN(n2874) );
  OAI22_X2 U551 ( .A1(n2876), .A2(n4646), .B1(n4641), .B2(n2877), .ZN(
        u1_fracta_s[41]) );
  AOI22_X2 U552 ( .A1(n4615), .A2(u1_adj_op_out_sft_41_), .B1(n4619), .B2(
        u6_N38), .ZN(n2876) );
  OAI22_X2 U553 ( .A1(n2878), .A2(n4646), .B1(n4641), .B2(n2879), .ZN(
        u1_fracta_s[40]) );
  AOI22_X2 U554 ( .A1(n4615), .A2(u1_adj_op_out_sft_40_), .B1(n4619), .B2(
        u6_N37), .ZN(n2878) );
  OAI22_X2 U555 ( .A1(n2880), .A2(n4646), .B1(n4641), .B2(n2881), .ZN(
        u1_fracta_s[3]) );
  AOI22_X2 U556 ( .A1(n4628), .A2(u1_adj_op_out_sft_3_), .B1(n4621), .B2(u6_N0), .ZN(n2880) );
  OAI22_X2 U557 ( .A1(n2882), .A2(n4646), .B1(n4641), .B2(n2883), .ZN(
        u1_fracta_s[39]) );
  AOI22_X2 U558 ( .A1(n4628), .A2(u1_adj_op_out_sft_39_), .B1(n4619), .B2(
        u6_N36), .ZN(n2882) );
  OAI22_X2 U559 ( .A1(n2884), .A2(n4646), .B1(n4641), .B2(n2885), .ZN(
        u1_fracta_s[38]) );
  AOI22_X2 U560 ( .A1(n4606), .A2(u1_adj_op_out_sft_38_), .B1(n4619), .B2(
        u6_N35), .ZN(n2884) );
  OAI22_X2 U561 ( .A1(n2886), .A2(n4646), .B1(n4641), .B2(n2887), .ZN(
        u1_fracta_s[37]) );
  AOI22_X2 U562 ( .A1(n4606), .A2(u1_adj_op_out_sft_37_), .B1(n4619), .B2(
        u6_N34), .ZN(n2886) );
  OAI22_X2 U563 ( .A1(n2888), .A2(n4646), .B1(n4641), .B2(n2889), .ZN(
        u1_fracta_s[36]) );
  AOI22_X2 U564 ( .A1(n4628), .A2(u1_adj_op_out_sft_36_), .B1(n4619), .B2(
        u6_N33), .ZN(n2888) );
  OAI22_X2 U565 ( .A1(n2890), .A2(n4646), .B1(n4641), .B2(n2891), .ZN(
        u1_fracta_s[35]) );
  AOI22_X2 U566 ( .A1(n4615), .A2(u1_adj_op_out_sft_35_), .B1(n4619), .B2(
        u6_N32), .ZN(n2890) );
  OAI22_X2 U567 ( .A1(n2892), .A2(n4647), .B1(n4641), .B2(n2893), .ZN(
        u1_fracta_s[34]) );
  AOI22_X2 U568 ( .A1(n4606), .A2(u1_adj_op_out_sft_34_), .B1(n4619), .B2(
        u6_N31), .ZN(n2892) );
  OAI22_X2 U569 ( .A1(n2894), .A2(n4647), .B1(n4641), .B2(n2895), .ZN(
        u1_fracta_s[33]) );
  AOI22_X2 U570 ( .A1(n4628), .A2(u1_adj_op_out_sft_33_), .B1(n4621), .B2(
        u6_N30), .ZN(n2894) );
  OAI22_X2 U571 ( .A1(n2896), .A2(n4647), .B1(n4641), .B2(n2897), .ZN(
        u1_fracta_s[32]) );
  AOI22_X2 U572 ( .A1(n4606), .A2(u1_adj_op_out_sft_32_), .B1(n4619), .B2(
        u6_N29), .ZN(n2896) );
  OAI22_X2 U573 ( .A1(n2898), .A2(n4647), .B1(n4642), .B2(n2899), .ZN(
        u1_fracta_s[31]) );
  AOI22_X2 U574 ( .A1(n4606), .A2(u1_adj_op_out_sft_31_), .B1(n4619), .B2(
        u6_N28), .ZN(n2898) );
  OAI22_X2 U575 ( .A1(n2900), .A2(n4647), .B1(n4642), .B2(n2901), .ZN(
        u1_fracta_s[30]) );
  AOI22_X2 U576 ( .A1(n4628), .A2(u1_adj_op_out_sft_30_), .B1(n4619), .B2(
        u6_N27), .ZN(n2900) );
  OAI22_X2 U577 ( .A1(n4643), .A2(n2902), .B1(n4649), .B2(n2903), .ZN(
        u1_fracta_s[2]) );
  NAND2_X2 U578 ( .A1(u1_adj_op_out_sft_2_), .A2(n4610), .ZN(n2902) );
  OAI22_X2 U579 ( .A1(n2904), .A2(n4647), .B1(n4642), .B2(n2905), .ZN(
        u1_fracta_s[29]) );
  AOI22_X2 U580 ( .A1(n4615), .A2(u1_adj_op_out_sft_29_), .B1(n4619), .B2(
        u6_N26), .ZN(n2904) );
  OAI22_X2 U581 ( .A1(n2906), .A2(n4647), .B1(n4638), .B2(n2907), .ZN(
        u1_fracta_s[28]) );
  AOI22_X2 U582 ( .A1(n4606), .A2(u1_adj_op_out_sft_28_), .B1(n4619), .B2(
        u6_N25), .ZN(n2906) );
  OAI22_X2 U583 ( .A1(n2908), .A2(n4645), .B1(n4638), .B2(n2909), .ZN(
        u1_fracta_s[27]) );
  AOI22_X2 U584 ( .A1(n4606), .A2(u1_adj_op_out_sft_27_), .B1(n4619), .B2(
        u6_N24), .ZN(n2908) );
  OAI22_X2 U585 ( .A1(n2910), .A2(n4647), .B1(n4649), .B2(n2911), .ZN(
        u1_fracta_s[26]) );
  AOI22_X2 U586 ( .A1(n4606), .A2(u1_adj_op_out_sft_26_), .B1(n4619), .B2(
        u6_N23), .ZN(n2910) );
  OAI22_X2 U587 ( .A1(n2912), .A2(n4647), .B1(n4649), .B2(n2913), .ZN(
        u1_fracta_s[25]) );
  AOI22_X2 U588 ( .A1(n4606), .A2(u1_adj_op_out_sft_25_), .B1(n4619), .B2(
        u6_N22), .ZN(n2912) );
  OAI22_X2 U589 ( .A1(n2914), .A2(n4647), .B1(n4642), .B2(n2915), .ZN(
        u1_fracta_s[24]) );
  AOI22_X2 U590 ( .A1(n4606), .A2(u1_adj_op_out_sft_24_), .B1(n4619), .B2(
        u6_N21), .ZN(n2914) );
  OAI22_X2 U591 ( .A1(n2916), .A2(n4647), .B1(n4638), .B2(n2917), .ZN(
        u1_fracta_s[23]) );
  AOI22_X2 U592 ( .A1(n4606), .A2(u1_adj_op_out_sft_23_), .B1(n4619), .B2(
        u6_N20), .ZN(n2916) );
  OAI22_X2 U593 ( .A1(n2918), .A2(n4647), .B1(n4642), .B2(n2919), .ZN(
        u1_fracta_s[22]) );
  AOI22_X2 U594 ( .A1(n4628), .A2(u1_adj_op_out_sft_22_), .B1(n4622), .B2(
        u6_N19), .ZN(n2918) );
  OAI22_X2 U595 ( .A1(n2920), .A2(n4647), .B1(n4642), .B2(n2921), .ZN(
        u1_fracta_s[21]) );
  AOI22_X2 U596 ( .A1(n4606), .A2(u1_adj_op_out_sft_21_), .B1(n4622), .B2(
        u6_N18), .ZN(n2920) );
  OAI22_X2 U597 ( .A1(n2922), .A2(n4647), .B1(n4642), .B2(n2923), .ZN(
        u1_fracta_s[20]) );
  AOI22_X2 U598 ( .A1(n4615), .A2(u1_adj_op_out_sft_20_), .B1(n4622), .B2(
        u6_N17), .ZN(n2922) );
  OAI22_X2 U599 ( .A1(n4643), .A2(n2924), .B1(n4642), .B2(n2925), .ZN(
        u1_fracta_s[1]) );
  NAND2_X2 U600 ( .A1(u1_adj_op_out_sft_1_), .A2(n4628), .ZN(n2924) );
  OAI22_X2 U601 ( .A1(n2926), .A2(n4647), .B1(n4642), .B2(n2927), .ZN(
        u1_fracta_s[19]) );
  AOI22_X2 U602 ( .A1(n4606), .A2(u1_adj_op_out_sft_19_), .B1(n4622), .B2(
        u6_N16), .ZN(n2926) );
  OAI22_X2 U603 ( .A1(n2928), .A2(n4647), .B1(n4642), .B2(n2929), .ZN(
        u1_fracta_s[18]) );
  AOI22_X2 U604 ( .A1(n4628), .A2(u1_adj_op_out_sft_18_), .B1(n4622), .B2(
        u6_N15), .ZN(n2928) );
  OAI22_X2 U605 ( .A1(n2930), .A2(n4647), .B1(n4642), .B2(n2931), .ZN(
        u1_fracta_s[17]) );
  AOI22_X2 U606 ( .A1(n4606), .A2(u1_adj_op_out_sft_17_), .B1(n4622), .B2(
        u6_N14), .ZN(n2930) );
  OAI22_X2 U607 ( .A1(n2932), .A2(n4647), .B1(n4642), .B2(n2933), .ZN(
        u1_fracta_s[16]) );
  AOI22_X2 U608 ( .A1(n4606), .A2(u1_adj_op_out_sft_16_), .B1(n4622), .B2(
        u6_N13), .ZN(n2932) );
  OAI22_X2 U609 ( .A1(n2934), .A2(n4647), .B1(n4642), .B2(n2935), .ZN(
        u1_fracta_s[15]) );
  AOI22_X2 U610 ( .A1(n4606), .A2(u1_adj_op_out_sft_15_), .B1(n4622), .B2(
        u6_N12), .ZN(n2934) );
  OAI22_X2 U611 ( .A1(n2936), .A2(n4647), .B1(n4642), .B2(n2937), .ZN(
        u1_fracta_s[14]) );
  AOI22_X2 U612 ( .A1(n4606), .A2(u1_adj_op_out_sft_14_), .B1(n4622), .B2(
        u6_N11), .ZN(n2936) );
  OAI22_X2 U613 ( .A1(n2938), .A2(n4651), .B1(n4642), .B2(n2939), .ZN(
        u1_fracta_s[13]) );
  AOI22_X2 U614 ( .A1(n4606), .A2(u1_adj_op_out_sft_13_), .B1(n4621), .B2(
        u6_N10), .ZN(n2938) );
  OAI22_X2 U615 ( .A1(n2940), .A2(n4651), .B1(n4642), .B2(n2941), .ZN(
        u1_fracta_s[12]) );
  AOI22_X2 U616 ( .A1(n4606), .A2(u1_adj_op_out_sft_12_), .B1(n4622), .B2(
        u6_N9), .ZN(n2940) );
  OAI22_X2 U617 ( .A1(n2942), .A2(n4651), .B1(n4649), .B2(n2943), .ZN(
        u1_fracta_s[11]) );
  AOI22_X2 U618 ( .A1(n4606), .A2(u1_adj_op_out_sft_11_), .B1(n4622), .B2(
        u6_N8), .ZN(n2942) );
  OAI22_X2 U619 ( .A1(n2944), .A2(n4645), .B1(n4649), .B2(n2945), .ZN(
        u1_fracta_s[10]) );
  AOI22_X2 U620 ( .A1(n4606), .A2(u1_adj_op_out_sft_10_), .B1(n4622), .B2(
        u6_N7), .ZN(n2944) );
  OAI22_X2 U621 ( .A1(n4643), .A2(n2946), .B1(n4649), .B2(n2947), .ZN(
        u1_fracta_s[0]) );
  NAND2_X2 U622 ( .A1(n4611), .A2(n2948), .ZN(n2946) );
  AOI22_X2 U623 ( .A1(n4622), .A2(u1_adj_op_out_sft_9_), .B1(fracta_mul[6]), 
        .B2(n4612), .ZN(n2837) );
  AOI22_X2 U624 ( .A1(n4622), .A2(u1_adj_op_out_sft_8_), .B1(n4615), .B2(
        fracta_mul[5]), .ZN(n2839) );
  AOI22_X2 U625 ( .A1(n4622), .A2(u1_adj_op_out_sft_7_), .B1(n4628), .B2(
        fracta_mul[4]), .ZN(n2841) );
  AOI22_X2 U626 ( .A1(n4622), .A2(u1_adj_op_out_sft_6_), .B1(n4628), .B2(
        fracta_mul[3]), .ZN(n2843) );
  AOI22_X2 U627 ( .A1(n4622), .A2(u1_adj_op_out_sft_5_), .B1(n4615), .B2(
        fracta_mul[2]), .ZN(n2845) );
  AOI22_X2 U628 ( .A1(n4621), .A2(u1_adj_op_out_sft_55_), .B1(n4602), .B2(
        n4612), .ZN(n2847) );
  AOI22_X2 U629 ( .A1(n4621), .A2(u1_adj_op_out_sft_54_), .B1(n4615), .B2(
        fracta_mul[51]), .ZN(n2849) );
  AOI22_X2 U630 ( .A1(n4621), .A2(u1_adj_op_out_sft_53_), .B1(n4606), .B2(
        fracta_mul[50]), .ZN(n2851) );
  AOI22_X2 U631 ( .A1(n4621), .A2(u1_adj_op_out_sft_52_), .B1(n4615), .B2(
        fracta_mul[49]), .ZN(n2853) );
  AOI22_X2 U632 ( .A1(n4621), .A2(u1_adj_op_out_sft_51_), .B1(n4615), .B2(
        fracta_mul[48]), .ZN(n2855) );
  AOI22_X2 U633 ( .A1(n4621), .A2(u1_adj_op_out_sft_50_), .B1(n4615), .B2(
        fracta_mul[47]), .ZN(n2857) );
  AOI22_X2 U634 ( .A1(n4621), .A2(u1_adj_op_out_sft_4_), .B1(n4628), .B2(
        fracta_mul[1]), .ZN(n2859) );
  AOI22_X2 U635 ( .A1(n4621), .A2(u1_adj_op_out_sft_49_), .B1(n4606), .B2(
        fracta_mul[46]), .ZN(n2861) );
  AOI22_X2 U636 ( .A1(n4621), .A2(u1_adj_op_out_sft_48_), .B1(n4615), .B2(
        fracta_mul[45]), .ZN(n2863) );
  AOI22_X2 U637 ( .A1(n4621), .A2(u1_adj_op_out_sft_47_), .B1(n4615), .B2(
        fracta_mul[44]), .ZN(n2865) );
  AOI22_X2 U638 ( .A1(n4621), .A2(u1_adj_op_out_sft_46_), .B1(n4615), .B2(
        fracta_mul[43]), .ZN(n2867) );
  AOI22_X2 U639 ( .A1(n4621), .A2(u1_adj_op_out_sft_45_), .B1(n4615), .B2(
        fracta_mul[42]), .ZN(n2869) );
  AOI22_X2 U640 ( .A1(n4621), .A2(u1_adj_op_out_sft_44_), .B1(n4615), .B2(
        fracta_mul[41]), .ZN(n2871) );
  AOI22_X2 U641 ( .A1(n4621), .A2(u1_adj_op_out_sft_43_), .B1(n4615), .B2(
        fracta_mul[40]), .ZN(n2873) );
  AOI22_X2 U642 ( .A1(n4621), .A2(u1_adj_op_out_sft_42_), .B1(n4615), .B2(
        fracta_mul[39]), .ZN(n2875) );
  AOI22_X2 U643 ( .A1(n4621), .A2(u1_adj_op_out_sft_41_), .B1(n4615), .B2(
        fracta_mul[38]), .ZN(n2877) );
  AOI22_X2 U644 ( .A1(n4621), .A2(u1_adj_op_out_sft_40_), .B1(n4615), .B2(
        fracta_mul[37]), .ZN(n2879) );
  AOI22_X2 U645 ( .A1(n4621), .A2(u1_adj_op_out_sft_3_), .B1(n4615), .B2(
        fracta_mul[0]), .ZN(n2881) );
  AOI22_X2 U646 ( .A1(n4619), .A2(u1_adj_op_out_sft_39_), .B1(n4606), .B2(
        fracta_mul[36]), .ZN(n2883) );
  AOI22_X2 U647 ( .A1(n4622), .A2(u1_adj_op_out_sft_38_), .B1(n4606), .B2(
        fracta_mul[35]), .ZN(n2885) );
  AOI22_X2 U648 ( .A1(n4621), .A2(u1_adj_op_out_sft_37_), .B1(n4606), .B2(
        fracta_mul[34]), .ZN(n2887) );
  AOI22_X2 U649 ( .A1(n4621), .A2(u1_adj_op_out_sft_36_), .B1(n4606), .B2(
        fracta_mul[33]), .ZN(n2889) );
  AOI22_X2 U650 ( .A1(n4621), .A2(u1_adj_op_out_sft_35_), .B1(n4606), .B2(
        fracta_mul[32]), .ZN(n2891) );
  AOI22_X2 U651 ( .A1(n4621), .A2(u1_adj_op_out_sft_34_), .B1(n4606), .B2(
        fracta_mul[31]), .ZN(n2893) );
  AOI22_X2 U652 ( .A1(n4621), .A2(u1_adj_op_out_sft_33_), .B1(n4606), .B2(
        fracta_mul[30]), .ZN(n2895) );
  AOI22_X2 U653 ( .A1(n4621), .A2(u1_adj_op_out_sft_32_), .B1(n4606), .B2(
        fracta_mul[29]), .ZN(n2897) );
  AOI22_X2 U654 ( .A1(n4621), .A2(u1_adj_op_out_sft_31_), .B1(n4611), .B2(
        fracta_mul[28]), .ZN(n2899) );
  AOI22_X2 U655 ( .A1(n4619), .A2(u1_adj_op_out_sft_30_), .B1(n4606), .B2(
        fracta_mul[27]), .ZN(n2901) );
  NAND2_X2 U656 ( .A1(u1_adj_op_out_sft_2_), .A2(n4626), .ZN(n2903) );
  AOI22_X2 U657 ( .A1(n4619), .A2(u1_adj_op_out_sft_29_), .B1(n4606), .B2(
        fracta_mul[26]), .ZN(n2905) );
  AOI22_X2 U658 ( .A1(n4619), .A2(u1_adj_op_out_sft_28_), .B1(n4611), .B2(
        fracta_mul[25]), .ZN(n2907) );
  AOI22_X2 U659 ( .A1(n4619), .A2(u1_adj_op_out_sft_27_), .B1(n4628), .B2(
        fracta_mul[24]), .ZN(n2909) );
  AOI22_X2 U660 ( .A1(n4619), .A2(u1_adj_op_out_sft_26_), .B1(n4611), .B2(
        fracta_mul[23]), .ZN(n2911) );
  AOI22_X2 U661 ( .A1(n4619), .A2(u1_adj_op_out_sft_25_), .B1(n4611), .B2(
        fracta_mul[22]), .ZN(n2913) );
  AOI22_X2 U662 ( .A1(n4619), .A2(u1_adj_op_out_sft_24_), .B1(n4611), .B2(
        fracta_mul[21]), .ZN(n2915) );
  AOI22_X2 U663 ( .A1(n4619), .A2(u1_adj_op_out_sft_23_), .B1(n4611), .B2(
        fracta_mul[20]), .ZN(n2917) );
  AOI22_X2 U664 ( .A1(n4619), .A2(u1_adj_op_out_sft_22_), .B1(n4611), .B2(
        fracta_mul[19]), .ZN(n2919) );
  AOI22_X2 U665 ( .A1(n4619), .A2(u1_adj_op_out_sft_21_), .B1(n4611), .B2(
        fracta_mul[18]), .ZN(n2921) );
  AOI22_X2 U666 ( .A1(n4619), .A2(u1_adj_op_out_sft_20_), .B1(n4611), .B2(
        fracta_mul[17]), .ZN(n2923) );
  NAND2_X2 U667 ( .A1(u1_adj_op_out_sft_1_), .A2(n4626), .ZN(n2925) );
  AOI22_X2 U668 ( .A1(n4619), .A2(u1_adj_op_out_sft_19_), .B1(n4615), .B2(
        fracta_mul[16]), .ZN(n2927) );
  AOI22_X2 U669 ( .A1(n4619), .A2(u1_adj_op_out_sft_18_), .B1(n4610), .B2(
        fracta_mul[15]), .ZN(n2929) );
  AOI22_X2 U670 ( .A1(n4619), .A2(u1_adj_op_out_sft_17_), .B1(n4610), .B2(
        fracta_mul[14]), .ZN(n2931) );
  AOI22_X2 U671 ( .A1(n4619), .A2(u1_adj_op_out_sft_16_), .B1(n4610), .B2(
        fracta_mul[13]), .ZN(n2933) );
  AOI22_X2 U672 ( .A1(n4621), .A2(u1_adj_op_out_sft_15_), .B1(n4610), .B2(
        fracta_mul[12]), .ZN(n2935) );
  AOI22_X2 U673 ( .A1(n4621), .A2(u1_adj_op_out_sft_14_), .B1(n4610), .B2(
        fracta_mul[11]), .ZN(n2937) );
  AOI22_X2 U674 ( .A1(n4621), .A2(u1_adj_op_out_sft_13_), .B1(n4610), .B2(
        fracta_mul[10]), .ZN(n2939) );
  AOI22_X2 U675 ( .A1(n4621), .A2(u1_adj_op_out_sft_12_), .B1(n4610), .B2(
        fracta_mul[9]), .ZN(n2941) );
  AOI22_X2 U676 ( .A1(n4621), .A2(u1_adj_op_out_sft_11_), .B1(n4610), .B2(
        fracta_mul[8]), .ZN(n2943) );
  AOI22_X2 U677 ( .A1(n4621), .A2(u1_adj_op_out_sft_10_), .B1(n4610), .B2(
        fracta_mul[7]), .ZN(n2945) );
  NAND2_X2 U678 ( .A1(n2948), .A2(n4626), .ZN(n2947) );
  OR3_X2 U679 ( .A1(u1_adj_op_out_sft_0_), .A2(n2949), .A3(n2950), .ZN(n2948)
         );
  AOI221_X2 U681 ( .B1(n6214), .B2(n2954), .C1(n6218), .C2(n2955), .A(n2956), 
        .ZN(n2952) );
  OAI22_X2 U682 ( .A1(n2957), .A2(n2958), .B1(n2959), .B2(n2960), .ZN(n2956)
         );
  AOI221_X2 U683 ( .B1(n6213), .B2(n2962), .C1(n6222), .C2(n2963), .A(n2964), 
        .ZN(n2951) );
  OAI22_X2 U684 ( .A1(n2965), .A2(n2966), .B1(n2967), .B2(n2968), .ZN(n2964)
         );
  OAI22_X2 U687 ( .A1(n2975), .A2(n2976), .B1(n2961), .B2(n2977), .ZN(n2974)
         );
  AOI22_X2 U688 ( .A1(n6216), .A2(n2978), .B1(n6220), .B2(n2979), .ZN(n2969)
         );
  OAI222_X2 U691 ( .A1(n2985), .A2(n2966), .B1(n2986), .B2(n2968), .C1(n2987), 
        .C2(n2980), .ZN(n2984) );
  OAI221_X2 U692 ( .B1(n2988), .B2(n2975), .C1(n2989), .C2(n2961), .A(n2990), 
        .ZN(n2983) );
  AOI22_X2 U693 ( .A1(n6216), .A2(n2991), .B1(n6220), .B2(n2992), .ZN(n2990)
         );
  OAI221_X2 U695 ( .B1(n2996), .B2(n2966), .C1(n2997), .C2(n2980), .A(n2998), 
        .ZN(n2994) );
  AOI22_X2 U696 ( .A1(n6220), .A2(n2999), .B1(n6212), .B2(n3000), .ZN(n2998)
         );
  NAND4_X2 U699 ( .A1(n6217), .A2(n6224), .A3(n6225), .A4(n3004), .ZN(n2980)
         );
  OAI221_X2 U701 ( .B1(n3005), .B2(n2961), .C1(n3006), .C2(n2960), .A(n3007), 
        .ZN(n2993) );
  AOI22_X2 U702 ( .A1(n3008), .A2(n3009), .B1(n6214), .B2(n3010), .ZN(n3007)
         );
  NAND2_X2 U703 ( .A1(n6217), .A2(n3011), .ZN(n2975) );
  NAND2_X2 U707 ( .A1(n2988), .A2(n3013), .ZN(n2954) );
  NAND2_X2 U709 ( .A1(n2977), .A2(n3014), .ZN(n3010) );
  NAND2_X2 U711 ( .A1(n2989), .A2(n3015), .ZN(n2955) );
  AND2_X2 U712 ( .A1(n3005), .A2(n3016), .ZN(n2989) );
  NAND2_X2 U715 ( .A1(n3011), .A2(n3003), .ZN(n2961) );
  NAND2_X2 U718 ( .A1(n2959), .A2(n3017), .ZN(n2978) );
  NAND2_X2 U720 ( .A1(n3006), .A2(n3018), .ZN(n2991) );
  NAND2_X2 U722 ( .A1(n2957), .A2(n3019), .ZN(n2979) );
  OR2_X2 U724 ( .A1(n2999), .A2(u1_adj_op_37_), .ZN(n2992) );
  OR2_X2 U725 ( .A1(n2972), .A2(u1_adj_op_36_), .ZN(n2999) );
  NAND2_X2 U726 ( .A1(n2967), .A2(n3020), .ZN(n2972) );
  AND2_X2 U727 ( .A1(n2986), .A2(n3021), .ZN(n2967) );
  OR2_X2 U729 ( .A1(n2973), .A2(u1_adj_op_32_), .ZN(n3000) );
  NAND2_X2 U730 ( .A1(n2965), .A2(n3022), .ZN(n2973) );
  AND2_X2 U731 ( .A1(n2985), .A2(n3023), .ZN(n2965) );
  AND2_X2 U732 ( .A1(n2996), .A2(n3024), .ZN(n2985) );
  OR2_X2 U734 ( .A1(n2962), .A2(u1_adj_op_27_), .ZN(n2971) );
  NAND2_X2 U735 ( .A1(n2987), .A2(n3025), .ZN(n2962) );
  AND2_X2 U736 ( .A1(n2997), .A2(n3026), .ZN(n2987) );
  AND4_X2 U737 ( .A1(n3027), .A2(n3028), .A3(n3029), .A4(n3030), .ZN(n2997) );
  NOR4_X2 U738 ( .A1(n3031), .A2(u1_adj_op_3_), .A3(n6233), .A4(n6235), .ZN(
        n3030) );
  NAND4_X2 U739 ( .A1(n3032), .A2(n3033), .A3(n3034), .A4(n3035), .ZN(n3031)
         );
  NOR4_X2 U740 ( .A1(n3036), .A2(u1_adj_op_20_), .A3(u1_adj_op_22_), .A4(
        u1_adj_op_21_), .ZN(n3029) );
  NOR4_X2 U742 ( .A1(n3040), .A2(u1_adj_op_15_), .A3(u1_adj_op_17_), .A4(
        u1_adj_op_16_), .ZN(n3028) );
  NOR4_X2 U744 ( .A1(n3044), .A2(u1_adj_op_0_), .A3(u1_adj_op_11_), .A4(
        u1_adj_op_10_), .ZN(n3027) );
  AOI22_X2 U746 ( .A1(n4606), .A2(opb_r[61]), .B1(n4623), .B2(opa_r[61]), .ZN(
        n3048) );
  AOI22_X2 U747 ( .A1(n4606), .A2(opb_r[60]), .B1(n4623), .B2(opa_r[60]), .ZN(
        n3049) );
  OAI22_X2 U748 ( .A1(n4625), .A2(n4340), .B1(n4614), .B2(n4442), .ZN(
        u1_exp_small[7]) );
  OAI22_X2 U749 ( .A1(n4624), .A2(n4399), .B1(n4613), .B2(n4454), .ZN(
        u1_exp_small[6]) );
  OAI22_X2 U750 ( .A1(n4625), .A2(n4296), .B1(n4613), .B2(n4453), .ZN(
        u1_exp_small[5]) );
  OAI22_X2 U751 ( .A1(n4624), .A2(n4359), .B1(n4613), .B2(n4456), .ZN(
        u1_exp_small[4]) );
  OAI22_X2 U752 ( .A1(n4625), .A2(n4321), .B1(n4614), .B2(n4358), .ZN(
        u1_exp_small[3]) );
  OAI22_X2 U753 ( .A1(n4624), .A2(n4457), .B1(n4613), .B2(n4451), .ZN(
        u1_exp_small[2]) );
  OAI22_X2 U754 ( .A1(n4625), .A2(n4275), .B1(n4614), .B2(n4450), .ZN(
        u1_exp_small[1]) );
  OAI22_X2 U755 ( .A1(n4363), .A2(n4626), .B1(n4614), .B2(n4458), .ZN(
        u1_exp_small[10]) );
  OAI22_X2 U756 ( .A1(n4625), .A2(n4270), .B1(n4614), .B2(n4449), .ZN(
        u1_exp_small[0]) );
  NAND2_X2 U760 ( .A1(u1_exp_diff_2_), .A2(n6223), .ZN(n3003) );
  NAND2_X2 U761 ( .A1(u1_exp_diff_1_), .A2(n6223), .ZN(n2953) );
  NAND2_X2 U762 ( .A1(u1_exp_diff_0_), .A2(n6223), .ZN(n2995) );
  AND2_X2 U763 ( .A1(u1_exp_diff2[9]), .A2(n3052), .ZN(u1_exp_diff_9_) );
  AND2_X2 U764 ( .A1(u1_exp_diff2[8]), .A2(n3052), .ZN(u1_exp_diff_8_) );
  AND2_X2 U765 ( .A1(u1_exp_diff2[7]), .A2(n3052), .ZN(u1_exp_diff_7_) );
  AND2_X2 U766 ( .A1(u1_exp_diff2[6]), .A2(n3052), .ZN(u1_exp_diff_6_) );
  AND2_X2 U767 ( .A1(u1_exp_diff2[5]), .A2(n3052), .ZN(u1_exp_diff_5_) );
  AND2_X2 U768 ( .A1(u1_exp_diff2[4]), .A2(n3052), .ZN(u1_exp_diff_4_) );
  AND2_X2 U769 ( .A1(u1_exp_diff2[3]), .A2(n3052), .ZN(u1_exp_diff_3_) );
  AND2_X2 U770 ( .A1(u1_exp_diff2[2]), .A2(n3052), .ZN(u1_exp_diff_2_) );
  AND2_X2 U771 ( .A1(u1_exp_diff2[1]), .A2(n3052), .ZN(u1_exp_diff_1_) );
  AND2_X2 U772 ( .A1(u1_exp_diff2[10]), .A2(n3052), .ZN(u1_exp_diff_10_) );
  AND2_X2 U773 ( .A1(u1_exp_diff2[0]), .A2(n3052), .ZN(u1_exp_diff_0_) );
  AOI22_X2 U775 ( .A1(n4606), .A2(u6_N9), .B1(n4623), .B2(fracta_mul[9]), .ZN(
        n3035) );
  AOI22_X2 U776 ( .A1(n4607), .A2(u6_N8), .B1(n4623), .B2(fracta_mul[8]), .ZN(
        n3034) );
  AOI22_X2 U777 ( .A1(n4607), .A2(u6_N7), .B1(n4623), .B2(fracta_mul[7]), .ZN(
        n3033) );
  AOI22_X2 U778 ( .A1(n4607), .A2(u6_N6), .B1(n4623), .B2(fracta_mul[6]), .ZN(
        n3032) );
  AOI22_X2 U779 ( .A1(n4607), .A2(u6_N5), .B1(n4623), .B2(fracta_mul[5]), .ZN(
        n3053) );
  OAI22_X2 U780 ( .A1(n4625), .A2(n4459), .B1(n4613), .B2(n4273), .ZN(
        u1_adj_op_51_) );
  AOI22_X2 U781 ( .A1(n4609), .A2(u6_N50), .B1(n4623), .B2(fracta_mul[50]), 
        .ZN(n3013) );
  AOI22_X2 U782 ( .A1(n4609), .A2(u6_N4), .B1(n4623), .B2(fracta_mul[4]), .ZN(
        n3054) );
  AOI22_X2 U783 ( .A1(n4609), .A2(u6_N49), .B1(n4623), .B2(fracta_mul[49]), 
        .ZN(n3055) );
  AOI22_X2 U784 ( .A1(n4609), .A2(u6_N48), .B1(n4623), .B2(fracta_mul[48]), 
        .ZN(n3014) );
  AOI22_X2 U785 ( .A1(n4609), .A2(u6_N47), .B1(n4624), .B2(fracta_mul[47]), 
        .ZN(n3056) );
  AOI22_X2 U786 ( .A1(n4609), .A2(u6_N46), .B1(n4623), .B2(fracta_mul[46]), 
        .ZN(n3015) );
  AOI22_X2 U787 ( .A1(n4609), .A2(u6_N45), .B1(n4624), .B2(fracta_mul[45]), 
        .ZN(n3016) );
  OAI22_X2 U788 ( .A1(n4625), .A2(n4468), .B1(n4613), .B2(n4277), .ZN(
        u1_adj_op_44_) );
  AOI22_X2 U789 ( .A1(n4609), .A2(u6_N43), .B1(n4624), .B2(fracta_mul[43]), 
        .ZN(n3017) );
  OAI22_X2 U790 ( .A1(n4625), .A2(n4467), .B1(n4613), .B2(n4286), .ZN(
        u1_adj_op_42_) );
  AOI22_X2 U791 ( .A1(n4609), .A2(u6_N41), .B1(n4623), .B2(fracta_mul[41]), 
        .ZN(n3018) );
  AOI22_X2 U792 ( .A1(n4609), .A2(u6_N40), .B1(n4623), .B2(fracta_mul[40]), 
        .ZN(n3057) );
  OAI22_X2 U793 ( .A1(n4624), .A2(n4463), .B1(n4612), .B2(n4360), .ZN(
        u1_adj_op_3_) );
  AOI22_X2 U794 ( .A1(n4608), .A2(u6_N39), .B1(n4623), .B2(fracta_mul[39]), 
        .ZN(n3019) );
  OAI22_X2 U795 ( .A1(n4625), .A2(n4465), .B1(n4612), .B2(n4284), .ZN(
        u1_adj_op_38_) );
  OAI22_X2 U796 ( .A1(n4625), .A2(n4471), .B1(n4613), .B2(n4272), .ZN(
        u1_adj_op_37_) );
  OAI22_X2 U797 ( .A1(n4625), .A2(n4470), .B1(n4613), .B2(n4276), .ZN(
        u1_adj_op_36_) );
  AOI22_X2 U798 ( .A1(n4608), .A2(u6_N35), .B1(n4623), .B2(fracta_mul[35]), 
        .ZN(n3020) );
  AOI22_X2 U799 ( .A1(n4608), .A2(u6_N34), .B1(n4624), .B2(fracta_mul[34]), 
        .ZN(n3021) );
  AOI22_X2 U800 ( .A1(n4608), .A2(u6_N33), .B1(n4623), .B2(fracta_mul[33]), 
        .ZN(n3058) );
  OAI22_X2 U801 ( .A1(n4625), .A2(n4464), .B1(n4613), .B2(n4287), .ZN(
        u1_adj_op_32_) );
  AOI22_X2 U802 ( .A1(n4608), .A2(u6_N31), .B1(n4623), .B2(fracta_mul[31]), 
        .ZN(n3022) );
  AOI22_X2 U803 ( .A1(n4608), .A2(u6_N30), .B1(n4624), .B2(fracta_mul[30]), 
        .ZN(n3023) );
  AOI22_X2 U804 ( .A1(n4608), .A2(u6_N2), .B1(n4623), .B2(fracta_mul[2]), .ZN(
        n3038) );
  AOI22_X2 U805 ( .A1(n4608), .A2(u6_N29), .B1(n4624), .B2(fracta_mul[29]), 
        .ZN(n3024) );
  OAI22_X2 U806 ( .A1(n4625), .A2(n4469), .B1(n4615), .B2(n4285), .ZN(
        u1_adj_op_28_) );
  OAI22_X2 U807 ( .A1(n4625), .A2(n4466), .B1(n4613), .B2(n4301), .ZN(
        u1_adj_op_27_) );
  AOI22_X2 U808 ( .A1(n4609), .A2(u6_N26), .B1(n4624), .B2(fracta_mul[26]), 
        .ZN(n3025) );
  AOI22_X2 U809 ( .A1(n4608), .A2(u6_N25), .B1(n4624), .B2(fracta_mul[25]), 
        .ZN(n3026) );
  AOI22_X2 U810 ( .A1(n4608), .A2(u6_N24), .B1(n4624), .B2(fracta_mul[24]), 
        .ZN(n3037) );
  AOI22_X2 U811 ( .A1(n4608), .A2(u6_N23), .B1(n4624), .B2(fracta_mul[23]), 
        .ZN(n3039) );
  OAI22_X2 U812 ( .A1(n4625), .A2(n4462), .B1(n4614), .B2(n4283), .ZN(
        u1_adj_op_22_) );
  OAI22_X2 U813 ( .A1(n4625), .A2(n4325), .B1(n4613), .B2(n4292), .ZN(
        u1_adj_op_21_) );
  OAI22_X2 U814 ( .A1(n4625), .A2(n4366), .B1(n4614), .B2(n4320), .ZN(
        u1_adj_op_20_) );
  AOI22_X2 U815 ( .A1(n4607), .A2(u6_N1), .B1(n4624), .B2(fracta_mul[1]), .ZN(
        n3042) );
  AOI22_X2 U816 ( .A1(n4607), .A2(u6_N19), .B1(n4624), .B2(fracta_mul[19]), 
        .ZN(n3041) );
  AOI22_X2 U817 ( .A1(n4607), .A2(u6_N18), .B1(n4624), .B2(fracta_mul[18]), 
        .ZN(n3043) );
  OAI22_X2 U818 ( .A1(n4625), .A2(n4461), .B1(n4614), .B2(n4319), .ZN(
        u1_adj_op_17_) );
  OAI22_X2 U819 ( .A1(n4625), .A2(n4324), .B1(n4614), .B2(n4362), .ZN(
        u1_adj_op_16_) );
  OAI22_X2 U820 ( .A1(n4625), .A2(n4365), .B1(n4615), .B2(n4318), .ZN(
        u1_adj_op_15_) );
  AOI22_X2 U821 ( .A1(n4607), .A2(u6_N14), .B1(n4624), .B2(fracta_mul[14]), 
        .ZN(n3046) );
  AOI22_X2 U822 ( .A1(n4607), .A2(u6_N13), .B1(n4624), .B2(fracta_mul[13]), 
        .ZN(n3045) );
  AOI22_X2 U823 ( .A1(n4607), .A2(u6_N12), .B1(n4624), .B2(fracta_mul[12]), 
        .ZN(n3047) );
  OAI22_X2 U824 ( .A1(n4626), .A2(n4460), .B1(n4614), .B2(n4361), .ZN(
        u1_adj_op_11_) );
  OAI22_X2 U825 ( .A1(n4626), .A2(n4323), .B1(n4614), .B2(n4300), .ZN(
        u1_adj_op_10_) );
  OAI22_X2 U826 ( .A1(n4626), .A2(n4364), .B1(n4615), .B2(n4322), .ZN(
        u1_adj_op_0_) );
  OAI22_X2 U828 ( .A1(n4612), .A2(n4363), .B1(n4458), .B2(n4626), .ZN(
        u1_exp_large_10_) );
  AOI22_X2 U830 ( .A1(n4622), .A2(opb_r[61]), .B1(n4610), .B2(opa_r[61]), .ZN(
        n3050) );
  AOI22_X2 U832 ( .A1(n4622), .A2(opb_r[60]), .B1(n4610), .B2(opa_r[60]), .ZN(
        n3051) );
  OAI22_X2 U834 ( .A1(n4611), .A2(n4340), .B1(n4626), .B2(n4442), .ZN(
        u1_exp_large_7_) );
  OAI22_X2 U836 ( .A1(n4612), .A2(n4399), .B1(n4626), .B2(n4454), .ZN(
        u1_exp_large_6_) );
  OAI22_X2 U838 ( .A1(n4611), .A2(n4296), .B1(n4626), .B2(n4453), .ZN(
        u1_exp_large_5_) );
  OAI22_X2 U840 ( .A1(n4612), .A2(n4359), .B1(n4626), .B2(n4456), .ZN(
        u1_exp_large_4_) );
  OAI22_X2 U842 ( .A1(n4612), .A2(n4321), .B1(n4626), .B2(n4358), .ZN(
        u1_exp_large_3_) );
  OAI22_X2 U844 ( .A1(n4612), .A2(n4457), .B1(n4626), .B2(n4451), .ZN(
        u1_exp_large_2_) );
  OAI22_X2 U846 ( .A1(n4612), .A2(n4275), .B1(n4626), .B2(n4450), .ZN(
        u1_exp_large_1_) );
  OAI22_X2 U848 ( .A1(n4612), .A2(n4270), .B1(n4626), .B2(n4449), .ZN(
        u1_exp_large_0_) );
  NAND2_X2 U850 ( .A1(u6_N52), .A2(n4602), .ZN(u1_N46) );
  XOR2_X2 U851 ( .A(n4481), .B(u2_sign_d), .Z(u1_N232) );
  XOR2_X2 U852 ( .A(opa_r[63]), .B(opb_r[63]), .Z(u2_sign_d) );
  AOI221_X2 U856 ( .B1(opb_nan), .B2(n3063), .C1(n3064), .C2(
        u1_fracta_lt_fractb), .A(u1_signa_r), .ZN(n3060) );
  NAND2_X2 U858 ( .A1(opa_nan), .A2(opb_nan), .ZN(n3063) );
  OAI22_X2 U859 ( .A1(n4490), .A2(n3065), .B1(n3066), .B2(n3067), .ZN(u1_N218)
         );
  XOR2_X2 U860 ( .A(u1_signb_r), .B(u1_add_r), .Z(n3067) );
  AND2_X2 U861 ( .A1(n3065), .A2(n4490), .ZN(n3066) );
  AOI22_X2 U862 ( .A1(u0_snan_r_a), .A2(u0_expa_ff), .B1(u0_snan_r_b), .B2(
        u0_expb_ff), .ZN(n3068) );
  AOI22_X2 U863 ( .A1(u0_qnan_r_a), .A2(u0_expa_ff), .B1(u0_qnan_r_b), .B2(
        u0_expb_ff), .ZN(n3069) );
  NAND2_X2 U864 ( .A1(n3070), .A2(n3071), .ZN(u0_N7) );
  AND2_X2 U866 ( .A1(n4459), .A2(n3072), .ZN(u0_N5) );
  AND2_X2 U868 ( .A1(u0_fractb_00), .A2(u0_expb_00), .ZN(u0_N17) );
  AND2_X2 U869 ( .A1(u0_fracta_00), .A2(u0_expa_00), .ZN(u0_N16) );
  NAND2_X2 U870 ( .A1(u0_infb_f_r), .A2(u0_expb_ff), .ZN(n3070) );
  NAND2_X2 U871 ( .A1(u0_infa_f_r), .A2(u0_expa_ff), .ZN(n3071) );
  NAND4_X2 U874 ( .A1(opb_r[52]), .A2(opb_r[53]), .A3(n3076), .A4(n3077), .ZN(
        n3074) );
  NOR4_X2 U875 ( .A1(n3078), .A2(n4296), .A3(n4340), .A4(n4399), .ZN(n3077) );
  NAND4_X2 U878 ( .A1(opa_r[52]), .A2(opa_r[53]), .A3(n3079), .A4(n3080), .ZN(
        n3075) );
  NOR4_X2 U879 ( .A1(n3081), .A2(n4453), .A3(n4442), .A4(n4454), .ZN(n3080) );
  OAI22_X2 U882 ( .A1(n6303), .A2(n4626), .B1(n4614), .B2(n4603), .ZN(n4266)
         );
  AND2_X2 U883 ( .A1(n3073), .A2(n4273), .ZN(n4267) );
  AND4_X2 U884 ( .A1(n3082), .A2(n3083), .A3(n3084), .A4(n3085), .ZN(n3073) );
  NOR4_X2 U885 ( .A1(n3086), .A2(n3087), .A3(fracta_mul[2]), .A4(
        fracta_mul[23]), .ZN(n3085) );
  NAND4_X2 U887 ( .A1(n4277), .A2(n4367), .A3(n4478), .A4(n3088), .ZN(n3086)
         );
  NOR4_X2 U889 ( .A1(n3089), .A2(fracta_mul[20]), .A3(fracta_mul[22]), .A4(
        fracta_mul[21]), .ZN(n3084) );
  NAND2_X2 U890 ( .A1(n4322), .A2(n4373), .ZN(n3089) );
  AND2_X2 U892 ( .A1(n3091), .A2(n3092), .ZN(n3082) );
  NAND4_X2 U893 ( .A1(n4270), .A2(n4275), .A3(n3093), .A4(n3094), .ZN(u6_N52)
         );
  NOR4_X2 U894 ( .A1(n3095), .A2(opb_r[60]), .A3(opb_r[62]), .A4(opb_r[61]), 
        .ZN(n3094) );
  NAND4_X2 U898 ( .A1(n3096), .A2(n3097), .A3(n3098), .A4(n3099), .ZN(n3072)
         );
  NOR4_X2 U899 ( .A1(n3100), .A2(n3101), .A3(n3102), .A4(n3103), .ZN(n3099) );
  NAND4_X2 U900 ( .A1(n4323), .A2(n4460), .A3(n4364), .A4(n3104), .ZN(n3103)
         );
  NAND4_X2 U902 ( .A1(n4324), .A2(n4461), .A3(n4365), .A4(n3105), .ZN(n3102)
         );
  NAND4_X2 U904 ( .A1(n4325), .A2(n4462), .A3(n4366), .A4(n3106), .ZN(n3101)
         );
  OR4_X2 U906 ( .A1(u6_N27), .A2(u6_N28), .A3(u6_N26), .A4(n3107), .ZN(n3100)
         );
  OR4_X2 U907 ( .A1(u6_N31), .A2(u6_N30), .A3(u6_N2), .A4(u6_N29), .ZN(n3107)
         );
  OR3_X2 U909 ( .A1(u6_N50), .A2(u6_N5), .A3(u6_N4), .ZN(n3110) );
  OR4_X2 U910 ( .A1(u6_N6), .A2(u6_N7), .A3(u6_N8), .A4(u6_N9), .ZN(n3109) );
  OR4_X2 U911 ( .A1(u6_N45), .A2(u6_N46), .A3(u6_N44), .A4(n3111), .ZN(n3108)
         );
  OR3_X2 U912 ( .A1(u6_N47), .A2(u6_N49), .A3(u6_N48), .ZN(n3111) );
  NOR4_X2 U913 ( .A1(n3112), .A2(u6_N38), .A3(u6_N3), .A4(u6_N39), .ZN(n3097)
         );
  OR4_X2 U914 ( .A1(u6_N40), .A2(u6_N41), .A3(u6_N42), .A4(u6_N43), .ZN(n3112)
         );
  NOR4_X2 U915 ( .A1(n3113), .A2(u6_N32), .A3(u6_N34), .A4(u6_N33), .ZN(n3096)
         );
  OR3_X2 U916 ( .A1(u6_N36), .A2(u6_N37), .A3(u6_N35), .ZN(n3113) );
  AOI22_X2 U917 ( .A1(u3_N69), .A2(n4659), .B1(u3_N12), .B2(n4657), .ZN(n3114)
         );
  AOI22_X2 U918 ( .A1(u3_N68), .A2(n4659), .B1(u3_N11), .B2(n4658), .ZN(n3115)
         );
  AOI22_X2 U919 ( .A1(u3_N67), .A2(n4659), .B1(u3_N10), .B2(n4657), .ZN(n3116)
         );
  AOI22_X2 U920 ( .A1(u3_N66), .A2(n4305), .B1(u3_N9), .B2(n4658), .ZN(n3117)
         );
  AOI22_X2 U921 ( .A1(u3_N65), .A2(n4659), .B1(u3_N8), .B2(n4657), .ZN(n3118)
         );
  AOI22_X2 U922 ( .A1(u3_N115), .A2(n4305), .B1(u3_N58), .B2(n4658), .ZN(n3119) );
  AOI22_X2 U923 ( .A1(u3_N114), .A2(n4659), .B1(u3_N57), .B2(n4657), .ZN(n3120) );
  AOI22_X2 U924 ( .A1(u3_N113), .A2(n4305), .B1(u3_N56), .B2(n4658), .ZN(n3121) );
  AOI22_X2 U925 ( .A1(u3_N112), .A2(n4659), .B1(u3_N55), .B2(n4657), .ZN(n3122) );
  AOI22_X2 U926 ( .A1(u3_N111), .A2(n4305), .B1(u3_N54), .B2(n4658), .ZN(n3123) );
  AOI22_X2 U927 ( .A1(u3_N110), .A2(n4659), .B1(u3_N53), .B2(n4657), .ZN(n3124) );
  AOI22_X2 U928 ( .A1(u3_N64), .A2(n4305), .B1(u3_N7), .B2(n4657), .ZN(n3125)
         );
  AOI22_X2 U929 ( .A1(u3_N109), .A2(n4659), .B1(u3_N52), .B2(n4657), .ZN(n3126) );
  AOI22_X2 U930 ( .A1(u3_N108), .A2(n4305), .B1(u3_N51), .B2(n4657), .ZN(n3127) );
  AOI22_X2 U931 ( .A1(u3_N107), .A2(n4659), .B1(u3_N50), .B2(n4657), .ZN(n3128) );
  AOI22_X2 U932 ( .A1(u3_N106), .A2(n4305), .B1(u3_N49), .B2(n4657), .ZN(n3129) );
  AOI22_X2 U933 ( .A1(u3_N105), .A2(n4659), .B1(u3_N48), .B2(n4657), .ZN(n3130) );
  AOI22_X2 U934 ( .A1(u3_N104), .A2(n4305), .B1(u3_N47), .B2(n4657), .ZN(n3131) );
  AOI22_X2 U935 ( .A1(u3_N103), .A2(n4305), .B1(u3_N46), .B2(n4657), .ZN(n3132) );
  AOI22_X2 U936 ( .A1(u3_N102), .A2(n4305), .B1(u3_N45), .B2(n4657), .ZN(n3133) );
  AOI22_X2 U937 ( .A1(u3_N101), .A2(n4305), .B1(u3_N44), .B2(n4657), .ZN(n3134) );
  AOI22_X2 U938 ( .A1(u3_N100), .A2(n4305), .B1(u3_N43), .B2(n4657), .ZN(n3135) );
  AOI22_X2 U939 ( .A1(u3_N63), .A2(n4305), .B1(u3_N6), .B2(n4658), .ZN(n3136)
         );
  AOI22_X2 U940 ( .A1(u3_N99), .A2(n4305), .B1(u3_N42), .B2(n4658), .ZN(n3137)
         );
  AOI22_X2 U941 ( .A1(u3_N98), .A2(n4305), .B1(u3_N41), .B2(n4658), .ZN(n3138)
         );
  AOI22_X2 U942 ( .A1(u3_N97), .A2(n4305), .B1(u3_N40), .B2(n4658), .ZN(n3139)
         );
  AOI22_X2 U943 ( .A1(u3_N96), .A2(n4305), .B1(u3_N39), .B2(n4658), .ZN(n3140)
         );
  AOI22_X2 U944 ( .A1(u3_N95), .A2(n4305), .B1(u3_N38), .B2(n4658), .ZN(n3141)
         );
  AOI22_X2 U945 ( .A1(u3_N94), .A2(n4305), .B1(u3_N37), .B2(n4658), .ZN(n3142)
         );
  AOI22_X2 U946 ( .A1(u3_N93), .A2(n4305), .B1(u3_N36), .B2(n4658), .ZN(n3143)
         );
  AOI22_X2 U947 ( .A1(u3_N92), .A2(n4305), .B1(u3_N35), .B2(n4658), .ZN(n3144)
         );
  AOI22_X2 U948 ( .A1(u3_N91), .A2(n4305), .B1(u3_N34), .B2(n4658), .ZN(n3145)
         );
  AOI22_X2 U949 ( .A1(u3_N90), .A2(n4305), .B1(u3_N33), .B2(n4658), .ZN(n3146)
         );
  AOI22_X2 U950 ( .A1(u3_N62), .A2(n4305), .B1(u3_N5), .B2(n4657), .ZN(n3147)
         );
  AOI22_X2 U951 ( .A1(u3_N89), .A2(n4305), .B1(u3_N32), .B2(n4658), .ZN(n3148)
         );
  AOI22_X2 U952 ( .A1(u3_N88), .A2(n4659), .B1(u3_N31), .B2(n4657), .ZN(n3149)
         );
  AOI22_X2 U953 ( .A1(u3_N87), .A2(n4659), .B1(u3_N30), .B2(n4658), .ZN(n3150)
         );
  AOI22_X2 U954 ( .A1(u3_N86), .A2(n4659), .B1(u3_N29), .B2(n4657), .ZN(n3151)
         );
  AOI22_X2 U955 ( .A1(u3_N85), .A2(n4659), .B1(u3_N28), .B2(n4658), .ZN(n3152)
         );
  AOI22_X2 U956 ( .A1(u3_N84), .A2(n4659), .B1(u3_N27), .B2(n4657), .ZN(n3153)
         );
  AOI22_X2 U957 ( .A1(u3_N83), .A2(n4659), .B1(u3_N26), .B2(n4658), .ZN(n3154)
         );
  AOI22_X2 U958 ( .A1(u3_N82), .A2(n4659), .B1(u3_N25), .B2(n4657), .ZN(n3155)
         );
  AOI22_X2 U959 ( .A1(u3_N81), .A2(n4659), .B1(u3_N24), .B2(n4658), .ZN(n3156)
         );
  AOI22_X2 U960 ( .A1(u3_N80), .A2(n4659), .B1(u3_N23), .B2(n4658), .ZN(n3157)
         );
  AOI22_X2 U961 ( .A1(u3_N61), .A2(n4659), .B1(u3_N4), .B2(fasu_op), .ZN(n3158) );
  AOI22_X2 U962 ( .A1(u3_N79), .A2(n4659), .B1(u3_N22), .B2(fasu_op), .ZN(
        n3159) );
  AOI22_X2 U963 ( .A1(u3_N78), .A2(n4659), .B1(u3_N21), .B2(fasu_op), .ZN(
        n3160) );
  AOI22_X2 U964 ( .A1(u3_N77), .A2(n4659), .B1(u3_N20), .B2(fasu_op), .ZN(
        n3161) );
  AOI22_X2 U965 ( .A1(u3_N76), .A2(n4659), .B1(u3_N19), .B2(fasu_op), .ZN(
        n3162) );
  AOI22_X2 U966 ( .A1(u3_N75), .A2(n4659), .B1(u3_N18), .B2(fasu_op), .ZN(
        n3163) );
  AOI22_X2 U967 ( .A1(u3_N74), .A2(n4659), .B1(u3_N17), .B2(fasu_op), .ZN(
        n3164) );
  AOI22_X2 U968 ( .A1(u3_N73), .A2(n4659), .B1(u3_N16), .B2(fasu_op), .ZN(
        n3165) );
  AOI22_X2 U969 ( .A1(u3_N72), .A2(n4659), .B1(u3_N15), .B2(fasu_op), .ZN(
        n3166) );
  AOI22_X2 U970 ( .A1(u3_N71), .A2(n4659), .B1(u3_N14), .B2(fasu_op), .ZN(
        n3167) );
  AOI22_X2 U971 ( .A1(u3_N70), .A2(n4659), .B1(u3_N13), .B2(fasu_op), .ZN(
        n3168) );
  AOI22_X2 U972 ( .A1(u3_N60), .A2(n4659), .B1(u3_N3), .B2(n4660), .ZN(n3169)
         );
  NAND2_X2 U974 ( .A1(quo[107]), .A2(opb_dn), .ZN(n3170) );
  OAI22_X2 U975 ( .A1(n4601), .A2(n4277), .B1(n4602), .B2(n5878), .ZN(u6_N99)
         );
  AOI22_X2 U976 ( .A1(n4602), .A2(fracta_mul[43]), .B1(n4603), .B2(N299), .ZN(
        n3181) );
  OAI22_X2 U977 ( .A1(n4601), .A2(n4286), .B1(n4602), .B2(n5879), .ZN(u6_N97)
         );
  OAI22_X2 U978 ( .A1(n4601), .A2(n4472), .B1(n4602), .B2(n5880), .ZN(u6_N96)
         );
  AOI22_X2 U979 ( .A1(n4602), .A2(fracta_mul[40]), .B1(n4603), .B2(N296), .ZN(
        n3182) );
  OAI22_X2 U980 ( .A1(n4601), .A2(n4478), .B1(n4602), .B2(n5881), .ZN(u6_N94)
         );
  OAI22_X2 U981 ( .A1(n4601), .A2(n4284), .B1(n4602), .B2(n5882), .ZN(u6_N93)
         );
  OAI22_X2 U982 ( .A1(n4601), .A2(n4272), .B1(n4602), .B2(n5883), .ZN(u6_N92)
         );
  OAI22_X2 U983 ( .A1(n4601), .A2(n4276), .B1(n4602), .B2(n5884), .ZN(u6_N91)
         );
  OAI22_X2 U984 ( .A1(n4601), .A2(n4474), .B1(n4602), .B2(n5885), .ZN(u6_N90)
         );
  AOI22_X2 U985 ( .A1(n4602), .A2(fracta_mul[34]), .B1(n4603), .B2(N290), .ZN(
        n3183) );
  AOI22_X2 U986 ( .A1(n4602), .A2(fracta_mul[33]), .B1(n4603), .B2(N289), .ZN(
        n3184) );
  OAI22_X2 U987 ( .A1(n4601), .A2(n4287), .B1(n4602), .B2(n5886), .ZN(u6_N87)
         );
  OAI22_X2 U988 ( .A1(n4601), .A2(n4370), .B1(n4602), .B2(n5887), .ZN(u6_N86)
         );
  OAI22_X2 U989 ( .A1(n4601), .A2(n4479), .B1(n4602), .B2(n5888), .ZN(u6_N85)
         );
  OAI22_X2 U990 ( .A1(n4601), .A2(n4475), .B1(n4602), .B2(n5889), .ZN(u6_N84)
         );
  OAI22_X2 U991 ( .A1(n4601), .A2(n4285), .B1(n4602), .B2(n5890), .ZN(u6_N83)
         );
  OAI22_X2 U992 ( .A1(n4601), .A2(n4301), .B1(n4602), .B2(n5891), .ZN(u6_N82)
         );
  AOI22_X2 U993 ( .A1(n4602), .A2(fracta_mul[26]), .B1(n4603), .B2(N282), .ZN(
        n3185) );
  OAI22_X2 U994 ( .A1(n4601), .A2(n4473), .B1(n4602), .B2(n5892), .ZN(u6_N80)
         );
  AOI22_X2 U995 ( .A1(n4602), .A2(fracta_mul[24]), .B1(n4603), .B2(N280), .ZN(
        n3186) );
  AOI22_X2 U996 ( .A1(n4602), .A2(fracta_mul[23]), .B1(n4603), .B2(N279), .ZN(
        n3187) );
  OAI22_X2 U997 ( .A1(n4603), .A2(n4283), .B1(n4602), .B2(n5893), .ZN(u6_N77)
         );
  OAI22_X2 U998 ( .A1(n4603), .A2(n4292), .B1(n4602), .B2(n5894), .ZN(u6_N76)
         );
  OAI22_X2 U999 ( .A1(n4603), .A2(n4320), .B1(n4602), .B2(n5895), .ZN(u6_N75)
         );
  AOI22_X2 U1000 ( .A1(n4602), .A2(fracta_mul[19]), .B1(n4603), .B2(N275), 
        .ZN(n3188) );
  OAI22_X2 U1001 ( .A1(n4601), .A2(n4369), .B1(n4602), .B2(n5896), .ZN(u6_N73)
         );
  OAI22_X2 U1002 ( .A1(n4601), .A2(n4319), .B1(n4602), .B2(n5897), .ZN(u6_N72)
         );
  OAI22_X2 U1003 ( .A1(n4601), .A2(n4362), .B1(n4602), .B2(n5898), .ZN(u6_N71)
         );
  OAI22_X2 U1004 ( .A1(n4601), .A2(n4318), .B1(n4602), .B2(n5899), .ZN(u6_N70)
         );
  OAI22_X2 U1005 ( .A1(n4601), .A2(n4372), .B1(n4602), .B2(n5900), .ZN(u6_N69)
         );
  AOI22_X2 U1006 ( .A1(n4602), .A2(fracta_mul[13]), .B1(n4603), .B2(N269), 
        .ZN(n3189) );
  OAI22_X2 U1007 ( .A1(n4601), .A2(n4374), .B1(n4602), .B2(n5901), .ZN(u6_N67)
         );
  OAI22_X2 U1008 ( .A1(n4601), .A2(n4361), .B1(n4602), .B2(n5902), .ZN(u6_N66)
         );
  OAI22_X2 U1009 ( .A1(n4601), .A2(n4300), .B1(n4602), .B2(n5903), .ZN(u6_N65)
         );
  OAI22_X2 U1010 ( .A1(n4601), .A2(n4368), .B1(n4602), .B2(n5904), .ZN(u6_N64)
         );
  OAI22_X2 U1011 ( .A1(n4601), .A2(n4326), .B1(n4602), .B2(n5905), .ZN(u6_N63)
         );
  OAI22_X2 U1012 ( .A1(n4601), .A2(n4376), .B1(n4602), .B2(n5906), .ZN(u6_N62)
         );
  OAI22_X2 U1013 ( .A1(n4601), .A2(n4375), .B1(n4602), .B2(n5907), .ZN(u6_N61)
         );
  OAI22_X2 U1014 ( .A1(n4601), .A2(n4371), .B1(n4602), .B2(n5908), .ZN(u6_N60)
         );
  AOI22_X2 U1015 ( .A1(n4602), .A2(fracta_mul[4]), .B1(n4603), .B2(N260), .ZN(
        n3190) );
  OAI22_X2 U1016 ( .A1(n4601), .A2(n4360), .B1(n4602), .B2(n5909), .ZN(u6_N58)
         );
  AOI22_X2 U1017 ( .A1(n4602), .A2(fracta_mul[2]), .B1(n4603), .B2(N258), .ZN(
        n3191) );
  OAI22_X2 U1018 ( .A1(n4601), .A2(n4373), .B1(n4602), .B2(n5910), .ZN(u6_N56)
         );
  OAI22_X2 U1019 ( .A1(n4601), .A2(n4322), .B1(n4602), .B2(n5911), .ZN(u6_N55)
         );
  OR2_X2 U1020 ( .A1(N308), .A2(n4602), .ZN(u6_N107) );
  OAI22_X2 U1021 ( .A1(n4601), .A2(n4273), .B1(n4602), .B2(n5874), .ZN(u6_N106) );
  OAI22_X2 U1022 ( .A1(n4601), .A2(n4480), .B1(n4602), .B2(n5875), .ZN(u6_N105) );
  AOI22_X2 U1023 ( .A1(n4602), .A2(fracta_mul[49]), .B1(n4603), .B2(N305), 
        .ZN(n3192) );
  AOI22_X2 U1024 ( .A1(n4602), .A2(fracta_mul[48]), .B1(n4603), .B2(N304), 
        .ZN(n3193) );
  AOI22_X2 U1025 ( .A1(n4602), .A2(fracta_mul[47]), .B1(n4603), .B2(N303), 
        .ZN(n3194) );
  OAI22_X2 U1026 ( .A1(n4601), .A2(n4477), .B1(n4602), .B2(n5876), .ZN(u6_N101) );
  OAI22_X2 U1027 ( .A1(n4601), .A2(n4367), .B1(n4602), .B2(n5877), .ZN(u6_N100) );
  NAND4_X2 U1028 ( .A1(n4449), .A2(n4450), .A3(n3195), .A4(n3196), .ZN(u2_N157) );
  NOR4_X2 U1029 ( .A1(n3197), .A2(opa_r[60]), .A3(opa_r[62]), .A4(opa_r[61]), 
        .ZN(n3196) );
  NAND4_X2 U1032 ( .A1(n6282), .A2(n3198), .A3(n6280), .A4(n3199), .ZN(
        div_opa_ldz_d[4]) );
  NOR4_X2 U1033 ( .A1(n6292), .A2(n3200), .A3(n3201), .A4(n3202), .ZN(n3199)
         );
  NAND4_X2 U1038 ( .A1(n3210), .A2(n3211), .A3(n3212), .A4(n3213), .ZN(
        div_opa_ldz_d[3]) );
  NOR4_X2 U1039 ( .A1(n3214), .A2(n3215), .A3(n6294), .A4(n3216), .ZN(n3213)
         );
  NOR4_X2 U1040 ( .A1(fracta_mul[29]), .A2(n3217), .A3(n4285), .A4(n6279), 
        .ZN(n3216) );
  OAI22_X2 U1042 ( .A1(n4301), .A2(n3220), .B1(n3221), .B2(n3204), .ZN(n3214)
         );
  NAND2_X2 U1047 ( .A1(n3231), .A2(n3232), .ZN(div_opa_ldz_d[2]) );
  NOR4_X2 U1048 ( .A1(n3233), .A2(n3234), .A3(n6285), .A4(n3235), .ZN(n3232)
         );
  NOR4_X2 U1049 ( .A1(fracta_mul[33]), .A2(n6298), .A3(n4287), .A4(n6279), 
        .ZN(n3235) );
  AND3_X2 U1050 ( .A1(fracta_mul[48]), .A2(n4273), .A3(n3237), .ZN(n3234) );
  OAI222_X2 U1053 ( .A1(fracta_mul[26]), .A2(n3228), .B1(n3243), .B2(n3218), 
        .C1(n3244), .C2(n3204), .ZN(n3241) );
  AOI221_X2 U1054 ( .B1(n3223), .B2(n3245), .C1(fracta_mul[14]), .C2(n3246), 
        .A(n3247), .ZN(n3244) );
  OR2_X2 U1055 ( .A1(fracta_mul[18]), .A2(fracta_mul[19]), .ZN(n3248) );
  OR4_X2 U1059 ( .A1(n3249), .A2(n3250), .A3(n3251), .A4(n3252), .ZN(
        div_opa_ldz_d[1]) );
  NAND4_X2 U1060 ( .A1(n3207), .A2(n3253), .A3(n3254), .A4(n3255), .ZN(n3252)
         );
  NOR4_X2 U1061 ( .A1(n3256), .A2(n6291), .A3(n3257), .A4(n3258), .ZN(n3255)
         );
  NAND4_X2 U1063 ( .A1(n3260), .A2(fracta_mul[30]), .A3(n3261), .A4(n4370), 
        .ZN(n3207) );
  OAI211_X2 U1064 ( .C1(fracta_mul[51]), .C2(n3237), .A(n3230), .B(n3210), 
        .ZN(n3251) );
  AND4_X2 U1065 ( .A1(n3238), .A2(n6289), .A3(n3236), .A4(n3262), .ZN(n3210)
         );
  NOR4_X2 U1066 ( .A1(n3263), .A2(n3264), .A3(n3265), .A4(n6286), .ZN(n3262)
         );
  NAND2_X2 U1068 ( .A1(n3269), .A2(fracta_mul[38]), .ZN(n3238) );
  NAND2_X2 U1070 ( .A1(n3271), .A2(fracta_mul[22]), .ZN(n3239) );
  NAND4_X2 U1074 ( .A1(n6277), .A2(n3211), .A3(n3276), .A4(n3277), .ZN(
        div_opa_ldz_d[0]) );
  NOR4_X2 U1075 ( .A1(n3278), .A2(n3270), .A3(fracta_mul[51]), .A4(n3263), 
        .ZN(n3277) );
  NAND2_X2 U1078 ( .A1(n6284), .A2(n4301), .ZN(n3272) );
  NAND4_X2 U1083 ( .A1(n3253), .A2(n3259), .A3(n3280), .A4(n3281), .ZN(n3209)
         );
  AOI22_X2 U1084 ( .A1(n6284), .A2(fracta_mul[27]), .B1(n3260), .B2(
        fracta_mul[35]), .ZN(n3281) );
  OR4_X2 U1087 ( .A1(n3204), .A2(n4373), .A3(n3090), .A4(fracta_mul[2]), .ZN(
        n3253) );
  NAND2_X2 U1088 ( .A1(n3282), .A2(n4360), .ZN(n3090) );
  AOI22_X2 U1090 ( .A1(fracta_mul[43]), .A2(n3226), .B1(fracta_mul[11]), .B2(
        n6287), .ZN(n3211) );
  NAND4_X2 U1091 ( .A1(n6278), .A2(n3198), .A3(n3285), .A4(n3286), .ZN(n3242)
         );
  NAND2_X2 U1094 ( .A1(n3267), .A2(n4375), .ZN(n3205) );
  OR3_X2 U1097 ( .A1(n3264), .A2(n3256), .A3(n6283), .ZN(n3287) );
  AND3_X2 U1104 ( .A1(fracta_mul[31]), .A2(n3261), .A3(n3260), .ZN(n3291) );
  AND3_X2 U1106 ( .A1(fracta_mul[21]), .A2(n4283), .A3(n3271), .ZN(n3265) );
  NAND2_X2 U1109 ( .A1(n6288), .A2(n3222), .ZN(n3284) );
  NOR4_X2 U1112 ( .A1(fracta_mul[16]), .A2(fracta_mul[17]), .A3(fracta_mul[18]), .A4(fracta_mul[19]), .ZN(n3246) );
  NAND2_X2 U1115 ( .A1(n3260), .A2(n3091), .ZN(n3220) );
  NAND2_X2 U1121 ( .A1(n3269), .A2(n4284), .ZN(n3206) );
  NOR4_X2 U1123 ( .A1(fracta_mul[24]), .A2(fracta_mul[25]), .A3(fracta_mul[26]), .A4(fracta_mul[27]), .ZN(n3289) );
  OR2_X2 U1125 ( .A1(fracta_mul[42]), .A2(fracta_mul[43]), .ZN(n3243) );
  OR3_X2 U1127 ( .A1(fracta_mul[46]), .A2(fracta_mul[47]), .A3(n6295), .ZN(
        n3219) );
  AOI22_X2 U1130 ( .A1(u3_N116), .A2(n4659), .B1(u3_N59), .B2(n4660), .ZN(
        n3292) );
  NOR4_X2 U1131 ( .A1(n3293), .A2(n3294), .A3(n4489), .A4(n4384), .ZN(N923) );
  NAND4_X2 U1133 ( .A1(exp_mul[3]), .A2(exp_mul[2]), .A3(exp_mul[4]), .A4(
        n3295), .ZN(n3293) );
  AND4_X2 U1135 ( .A1(opb_00), .A2(opa_nan_r), .A3(n4486), .A4(n4382), .ZN(
        N913) );
  OAI211_X2 U1137 ( .C1(n3297), .C2(n3298), .A(n3299), .B(n3300), .ZN(N911) );
  NOR4_X2 U1139 ( .A1(n3304), .A2(n3305), .A3(n2507), .A4(n3306), .ZN(n3301)
         );
  OR2_X2 U1140 ( .A1(inf_mul2), .A2(inf_mul_r), .ZN(n3305) );
  NAND4_X2 U1141 ( .A1(n6341), .A2(n3307), .A3(n3308), .A4(n3309), .ZN(n3299)
         );
  OAI221_X2 U1143 ( .B1(n3310), .B2(n3311), .C1(n3312), .C2(n6458), .A(n3313), 
        .ZN(N906) );
  AND3_X2 U1146 ( .A1(fasu_op_r2), .A2(n3315), .A3(inf_d), .ZN(n3317) );
  NAND4_X2 U1148 ( .A1(n3321), .A2(n3322), .A3(n3323), .A4(n3324), .ZN(n3318)
         );
  NOR4_X2 U1149 ( .A1(n3325), .A2(n3326), .A3(n3327), .A4(n3328), .ZN(n3324)
         );
  NAND4_X2 U1150 ( .A1(n3329), .A2(n3330), .A3(n3331), .A4(n3332), .ZN(n3325)
         );
  NOR4_X2 U1151 ( .A1(n3333), .A2(n3334), .A3(n3335), .A4(n3336), .ZN(n3323)
         );
  NAND4_X2 U1152 ( .A1(n3337), .A2(n3338), .A3(n3339), .A4(n3340), .ZN(n3333)
         );
  AOI22_X2 U1153 ( .A1(opb_00), .A2(n4486), .B1(opa_inf), .B2(n4327), .ZN(
        n3310) );
  AOI221_X2 U1155 ( .B1(underflow_fmul_r[2]), .B2(n3345), .C1(
        underflow_fmul_r[1]), .C2(n3346), .A(n3347), .ZN(n3344) );
  OR2_X2 U1156 ( .A1(underflow_fmul_r[0]), .A2(n3348), .ZN(n3347) );
  NOR4_X2 U1157 ( .A1(n6447), .A2(n3304), .A3(n3349), .A4(n4485), .ZN(n3348)
         );
  NOR4_X2 U1158 ( .A1(n3350), .A2(n3351), .A3(n3352), .A4(n3353), .ZN(n3349)
         );
  NAND4_X2 U1159 ( .A1(n3354), .A2(n3355), .A3(n3356), .A4(n3357), .ZN(n3353)
         );
  NOR4_X2 U1160 ( .A1(n3358), .A2(prod[21]), .A3(prod[23]), .A4(prod[22]), 
        .ZN(n3357) );
  OR4_X2 U1161 ( .A1(prod[24]), .A2(prod[25]), .A3(prod[26]), .A4(prod[27]), 
        .ZN(n3358) );
  NOR4_X2 U1162 ( .A1(n3359), .A2(prod[16]), .A3(prod[18]), .A4(prod[17]), 
        .ZN(n3356) );
  OR3_X2 U1163 ( .A1(prod[1]), .A2(prod[20]), .A3(prod[19]), .ZN(n3359) );
  NOR4_X2 U1164 ( .A1(n3360), .A2(prod[105]), .A3(prod[11]), .A4(prod[10]), 
        .ZN(n3355) );
  OR4_X2 U1165 ( .A1(prod[12]), .A2(prod[13]), .A3(prod[14]), .A4(prod[15]), 
        .ZN(n3360) );
  NOR4_X2 U1166 ( .A1(n3361), .A2(prod[0]), .A3(prod[101]), .A4(prod[100]), 
        .ZN(n3354) );
  NAND4_X2 U1168 ( .A1(n3362), .A2(n3363), .A3(n3364), .A4(n3365), .ZN(n3352)
         );
  NOR4_X2 U1169 ( .A1(n3366), .A2(prod[46]), .A3(prod[48]), .A4(prod[47]), 
        .ZN(n3365) );
  OR4_X2 U1170 ( .A1(prod[49]), .A2(prod[4]), .A3(prod[50]), .A4(prod[51]), 
        .ZN(n3366) );
  NOR4_X2 U1171 ( .A1(n3367), .A2(prod[3]), .A3(prod[41]), .A4(prod[40]), .ZN(
        n3364) );
  OR4_X2 U1172 ( .A1(prod[42]), .A2(prod[43]), .A3(prod[44]), .A4(prod[45]), 
        .ZN(n3367) );
  NOR4_X2 U1173 ( .A1(n3368), .A2(prod[33]), .A3(prod[35]), .A4(prod[34]), 
        .ZN(n3363) );
  OR4_X2 U1174 ( .A1(prod[36]), .A2(prod[37]), .A3(prod[38]), .A4(prod[39]), 
        .ZN(n3368) );
  NOR4_X2 U1175 ( .A1(n3369), .A2(prod[28]), .A3(prod[2]), .A4(prod[29]), .ZN(
        n3362) );
  OR3_X2 U1176 ( .A1(prod[31]), .A2(prod[32]), .A3(prod[30]), .ZN(n3369) );
  NAND4_X2 U1177 ( .A1(n3370), .A2(n3371), .A3(n3372), .A4(n3373), .ZN(n3351)
         );
  NOR4_X2 U1178 ( .A1(n3374), .A2(prod[6]), .A3(prod[71]), .A4(prod[70]), .ZN(
        n3373) );
  NAND4_X2 U1179 ( .A1(n4313), .A2(n4407), .A3(n4298), .A4(n4343), .ZN(n3374)
         );
  NOR4_X2 U1180 ( .A1(n3375), .A2(prod[64]), .A3(prod[66]), .A4(prod[65]), 
        .ZN(n3372) );
  NOR4_X2 U1182 ( .A1(n3376), .A2(prod[58]), .A3(prod[5]), .A4(prod[59]), .ZN(
        n3371) );
  NAND4_X2 U1183 ( .A1(n4346), .A2(n4406), .A3(n4312), .A4(n4297), .ZN(n3376)
         );
  NOR4_X2 U1184 ( .A1(n3377), .A2(prod[52]), .A3(prod[54]), .A4(prod[53]), 
        .ZN(n3370) );
  NAND4_X2 U1186 ( .A1(n3378), .A2(n3379), .A3(n3380), .A4(n3381), .ZN(n3350)
         );
  NOR4_X2 U1187 ( .A1(n3382), .A2(prod[94]), .A3(prod[96]), .A4(prod[95]), 
        .ZN(n3381) );
  OR4_X2 U1188 ( .A1(prod[97]), .A2(prod[98]), .A3(prod[99]), .A4(prod[9]), 
        .ZN(n3382) );
  NOR4_X2 U1189 ( .A1(n3383), .A2(prod[88]), .A3(prod[8]), .A4(prod[89]), .ZN(
        n3380) );
  NAND4_X2 U1190 ( .A1(n4345), .A2(n4405), .A3(n4308), .A4(n4295), .ZN(n3383)
         );
  NOR4_X2 U1191 ( .A1(n3384), .A2(prod[81]), .A3(prod[83]), .A4(prod[82]), 
        .ZN(n3379) );
  NAND4_X2 U1192 ( .A1(n4344), .A2(n4404), .A3(n4307), .A4(n4294), .ZN(n3384)
         );
  NOR4_X2 U1193 ( .A1(n3385), .A2(prod[76]), .A3(prod[78]), .A4(prod[77]), 
        .ZN(n3378) );
  OR3_X2 U1194 ( .A1(prod[7]), .A2(prod[80]), .A3(prod[79]), .ZN(n3385) );
  NAND4_X2 U1196 ( .A1(n3388), .A2(n3389), .A3(n3390), .A4(n3391), .ZN(n3387)
         );
  NOR4_X2 U1197 ( .A1(n3392), .A2(n3393), .A3(n3394), .A4(n3395), .ZN(n3391)
         );
  AND3_X2 U1198 ( .A1(n3396), .A2(n3397), .A3(n3398), .ZN(n3390) );
  NAND4_X2 U1199 ( .A1(n3399), .A2(n3400), .A3(n3401), .A4(n3402), .ZN(n3319)
         );
  NOR4_X2 U1200 ( .A1(n3403), .A2(n3404), .A3(n3405), .A4(n3406), .ZN(n3402)
         );
  NAND4_X2 U1201 ( .A1(n3407), .A2(n3408), .A3(n3409), .A4(n3410), .ZN(n3403)
         );
  NOR4_X2 U1202 ( .A1(n3411), .A2(n3412), .A3(n3413), .A4(n3414), .ZN(n3401)
         );
  NOR4_X2 U1204 ( .A1(n3418), .A2(n3419), .A3(n3420), .A4(n3421), .ZN(n3400)
         );
  NAND4_X2 U1205 ( .A1(n3422), .A2(n3423), .A3(n3424), .A4(n3425), .ZN(n3418)
         );
  NOR4_X2 U1206 ( .A1(n3426), .A2(n3427), .A3(n3428), .A4(n3429), .ZN(n3399)
         );
  NAND4_X2 U1208 ( .A1(n3321), .A2(n3322), .A3(n3433), .A4(n3434), .ZN(n3386)
         );
  NOR4_X2 U1209 ( .A1(n3435), .A2(n3436), .A3(n3328), .A4(n3326), .ZN(n3434)
         );
  NAND4_X2 U1210 ( .A1(n3437), .A2(n3329), .A3(n3330), .A4(n3331), .ZN(n3435)
         );
  NOR4_X2 U1211 ( .A1(n3438), .A2(n3334), .A3(n3335), .A4(n3336), .ZN(n3433)
         );
  NOR4_X2 U1213 ( .A1(n3439), .A2(n3440), .A3(n3441), .A4(n3442), .ZN(n3322)
         );
  NAND4_X2 U1214 ( .A1(n3443), .A2(n3444), .A3(n3445), .A4(n3446), .ZN(n3439)
         );
  NOR4_X2 U1215 ( .A1(n3447), .A2(n3448), .A3(n3449), .A4(n3450), .ZN(n3321)
         );
  OAI221_X2 U1218 ( .B1(n3460), .B2(n6449), .C1(n3461), .C2(n4291), .A(n3462), 
        .ZN(N889) );
  AOI22_X2 U1221 ( .A1(n3464), .A2(n6316), .B1(n4540), .B2(n3463), .ZN(n3460)
         );
  AND2_X2 U1223 ( .A1(n3320), .A2(n3304), .ZN(n3466) );
  NAND2_X2 U1226 ( .A1(n4327), .A2(n4382), .ZN(n3306) );
  INV_X4 U1229 ( .A(n3346), .ZN(n3342) );
  NAND2_X2 U1231 ( .A1(n6316), .A2(n3472), .ZN(n3471) );
  NOR4_X2 U1232 ( .A1(exp_ovf_r[1]), .A2(n6465), .A3(u4_exp_in_mi1_11_), .A4(
        n3476), .ZN(n3474) );
  OR3_X2 U1233 ( .A1(n4355), .A2(n3477), .A3(n3478), .ZN(n3470) );
  OAI211_X2 U1234 ( .C1(n3479), .C2(n3480), .A(n3481), .B(n3482), .ZN(n3469)
         );
  AOI221_X2 U1239 ( .B1(u4_N6279), .B2(n3490), .C1(n3491), .C2(exp_ovf_r[1]), 
        .A(n3492), .ZN(n3483) );
  INV_X4 U1240 ( .A(n3493), .ZN(n3492) );
  AND4_X2 U1242 ( .A1(u4_N6286), .A2(n3496), .A3(n3497), .A4(n3498), .ZN(n3494) );
  NOR4_X2 U1243 ( .A1(n3499), .A2(exp_r[3]), .A3(n4290), .A4(n4282), .ZN(n3498) );
  OR3_X2 U1244 ( .A1(n4281), .A2(n4353), .A3(exp_r[6]), .ZN(n3499) );
  INV_X4 U1246 ( .A(n2518), .ZN(n3496) );
  XOR2_X2 U1249 ( .A(n4656), .B(n5864), .Z(n3503) );
  NOR4_X2 U1250 ( .A1(n3505), .A2(n5868), .A3(n5870), .A4(n5869), .ZN(n3502)
         );
  NAND2_X2 U1252 ( .A1(u4_div_exp3[5]), .A2(n2394), .ZN(n3508) );
  NAND2_X2 U1255 ( .A1(u4_div_exp3[4]), .A2(n2394), .ZN(n3511) );
  NAND2_X2 U1258 ( .A1(u4_div_exp3[6]), .A2(n4542), .ZN(n3514) );
  NAND2_X2 U1262 ( .A1(u4_div_exp3[3]), .A2(n2394), .ZN(n3516) );
  NAND2_X2 U1265 ( .A1(u4_div_exp3[1]), .A2(n2394), .ZN(n3518) );
  NAND2_X2 U1268 ( .A1(u4_div_exp3[2]), .A2(n2394), .ZN(n3520) );
  NOR4_X2 U1270 ( .A1(n3504), .A2(n3521), .A3(n2430), .A4(n2427), .ZN(n3501)
         );
  NAND2_X2 U1272 ( .A1(u4_div_exp3[8]), .A2(n2394), .ZN(n3523) );
  NAND2_X2 U1275 ( .A1(u4_div_exp3[9]), .A2(n4542), .ZN(n3525) );
  NAND2_X2 U1277 ( .A1(n6465), .A2(n2423), .ZN(n3521) );
  NAND2_X2 U1279 ( .A1(u4_div_exp3[7]), .A2(n4542), .ZN(n3527) );
  NAND2_X2 U1282 ( .A1(u4_div_exp3[10]), .A2(n2394), .ZN(n3529) );
  OAI22_X2 U1287 ( .A1(exp_ovf_r[1]), .A2(n3530), .B1(n4452), .B2(n3531), .ZN(
        n3490) );
  AND2_X2 U1289 ( .A1(u4_N6280), .A2(n3495), .ZN(n3532) );
  INV_X4 U1290 ( .A(n3533), .ZN(n3530) );
  NAND4_X2 U1291 ( .A1(n3397), .A2(n3534), .A3(n3535), .A4(n3536), .ZN(n3480)
         );
  NAND4_X2 U1292 ( .A1(n3537), .A2(n3392), .A3(n3538), .A4(n3393), .ZN(n3479)
         );
  INV_X4 U1294 ( .A(n3541), .ZN(n3461) );
  OAI221_X2 U1295 ( .B1(n2433), .B2(n3475), .C1(n3542), .C2(n2434), .A(n3543), 
        .ZN(n3541) );
  AOI221_X2 U1296 ( .B1(n3544), .B2(n3545), .C1(n4540), .C2(n3495), .A(n3477), 
        .ZN(n3543) );
  NOR4_X2 U1299 ( .A1(n4656), .A2(n6307), .A3(n4441), .A4(n4351), .ZN(n3546)
         );
  INV_X4 U1300 ( .A(n3485), .ZN(n3475) );
  AOI22_X2 U1301 ( .A1(n3549), .A2(n4540), .B1(n4355), .B2(n3550), .ZN(n3456)
         );
  OAI211_X2 U1303 ( .C1(n3551), .C2(n4356), .A(n3553), .B(n3554), .ZN(n3549)
         );
  AND3_X2 U1305 ( .A1(n4352), .A2(n3488), .A3(n3557), .ZN(n3555) );
  NAND4_X2 U1307 ( .A1(n3302), .A2(n3303), .A3(opas_r2), .A4(n6308), .ZN(n3559) );
  AOI22_X2 U1308 ( .A1(n6314), .A2(n3560), .B1(n3561), .B2(n3343), .ZN(n3558)
         );
  OAI22_X2 U1309 ( .A1(n6341), .A2(n3562), .B1(n3563), .B2(n3311), .ZN(n3561)
         );
  AOI22_X2 U1310 ( .A1(n3564), .A2(n6455), .B1(n3565), .B2(n4491), .ZN(n3563)
         );
  NAND2_X2 U1312 ( .A1(opb_inf), .A2(opa_inf), .ZN(n3309) );
  NAND2_X2 U1313 ( .A1(n4491), .A2(n3308), .ZN(n3564) );
  AOI22_X2 U1314 ( .A1(n3314), .A2(n3566), .B1(nan_sign_d), .B2(n6457), .ZN(
        n3562) );
  INV_X4 U1315 ( .A(n3567), .ZN(n3566) );
  AOI22_X2 U1316 ( .A1(sign_fasu_r), .A2(n3298), .B1(result_zero_sign_d), .B2(
        n3568), .ZN(n3567) );
  INV_X4 U1317 ( .A(n3568), .ZN(n3298) );
  NAND2_X2 U1321 ( .A1(n3303), .A2(n4540), .ZN(n3311) );
  XOR2_X2 U1322 ( .A(sign_mul_r), .B(n3569), .Z(n3560) );
  NAND2_X2 U1324 ( .A1(n3303), .A2(n6316), .ZN(n3343) );
  NAND4_X2 U1326 ( .A1(n3570), .A2(n3571), .A3(n3572), .A4(n3573), .ZN(n3304)
         );
  NOR4_X2 U1327 ( .A1(n3574), .A2(n3575), .A3(n3576), .A4(n3577), .ZN(n3573)
         );
  NAND4_X2 U1328 ( .A1(n3445), .A2(n3446), .A3(n3578), .A4(n3579), .ZN(n3577)
         );
  NAND4_X2 U1329 ( .A1(n3580), .A2(n3337), .A3(n3338), .A4(n3339), .ZN(n3576)
         );
  NAND4_X2 U1330 ( .A1(n3340), .A2(n3581), .A3(n3582), .A4(n3437), .ZN(n3575)
         );
  NAND4_X2 U1331 ( .A1(n3329), .A2(n3330), .A3(n3331), .A4(n3397), .ZN(n3574)
         );
  NOR4_X2 U1333 ( .A1(n3586), .A2(n3587), .A3(n3588), .A4(n3589), .ZN(n3572)
         );
  NAND4_X2 U1335 ( .A1(n3410), .A2(n3590), .A3(n3591), .A4(n3592), .ZN(n3588)
         );
  NAND4_X2 U1336 ( .A1(n3453), .A2(n3451), .A3(n3452), .A4(n3593), .ZN(n3587)
         );
  NAND4_X2 U1337 ( .A1(n3594), .A2(n3595), .A3(n3443), .A4(n3444), .ZN(n3586)
         );
  NOR4_X2 U1338 ( .A1(n3596), .A2(n3597), .A3(n3598), .A4(n3599), .ZN(n3571)
         );
  NAND4_X2 U1340 ( .A1(n3423), .A2(n3424), .A3(n3425), .A4(n3602), .ZN(n3598)
         );
  NAND4_X2 U1341 ( .A1(n3603), .A2(n3604), .A3(n3417), .A4(n3415), .ZN(n3597)
         );
  NAND4_X2 U1342 ( .A1(n3416), .A2(n3605), .A3(n3606), .A4(n3607), .ZN(n3596)
         );
  NAND4_X2 U1344 ( .A1(n3398), .A2(n3611), .A3(n3612), .A4(n3613), .ZN(n3610)
         );
  NAND4_X2 U1345 ( .A1(n3432), .A2(n3430), .A3(n3431), .A4(n3614), .ZN(n3609)
         );
  NAND4_X2 U1346 ( .A1(n3540), .A2(n3615), .A3(n3539), .A4(n3616), .ZN(n3608)
         );
  NOR4_X2 U1347 ( .A1(n3535), .A2(n3536), .A3(n3537), .A4(n3392), .ZN(n3616)
         );
  INV_X4 U1348 ( .A(n3617), .ZN(n3392) );
  INV_X4 U1349 ( .A(n3388), .ZN(n3537) );
  INV_X4 U1350 ( .A(n3389), .ZN(n3536) );
  INV_X4 U1351 ( .A(n3396), .ZN(n3535) );
  NAND2_X2 U1352 ( .A1(n3618), .A2(n3619), .ZN(N855) );
  OR2_X2 U1353 ( .A1(n3583), .A2(n6310), .ZN(N854) );
  OR2_X2 U1354 ( .A1(n3584), .A2(n6310), .ZN(N853) );
  NAND2_X2 U1355 ( .A1(n3539), .A2(n3619), .ZN(N852) );
  NAND2_X2 U1356 ( .A1(n3540), .A2(n3619), .ZN(N851) );
  NAND2_X2 U1357 ( .A1(n3615), .A2(n3619), .ZN(N850) );
  NAND2_X2 U1358 ( .A1(n3617), .A2(n3619), .ZN(N849) );
  NAND2_X2 U1359 ( .A1(n3388), .A2(n3619), .ZN(N848) );
  NAND2_X2 U1360 ( .A1(n3389), .A2(n3619), .ZN(N847) );
  NAND2_X2 U1361 ( .A1(n3396), .A2(n3619), .ZN(N846) );
  NAND2_X2 U1362 ( .A1(n3398), .A2(n3619), .ZN(N845) );
  INV_X4 U1364 ( .A(n3427), .ZN(n3611) );
  OAI221_X2 U1365 ( .B1(n4593), .B2(n3621), .C1(n2520), .C2(n4591), .A(n4588), 
        .ZN(n3427) );
  INV_X4 U1366 ( .A(u4_fract_out_pl1_51_), .ZN(n3621) );
  INV_X4 U1368 ( .A(n3429), .ZN(n3612) );
  OAI221_X2 U1369 ( .B1(n4593), .B2(n3624), .C1(n2521), .C2(n4591), .A(n4588), 
        .ZN(n3429) );
  INV_X4 U1370 ( .A(u4_fract_out_pl1_50_), .ZN(n3624) );
  INV_X4 U1372 ( .A(n3428), .ZN(n3613) );
  OAI221_X2 U1373 ( .B1(n4593), .B2(n3625), .C1(n3626), .C2(n4591), .A(n4588), 
        .ZN(n3428) );
  INV_X4 U1374 ( .A(u4_fract_out_pl1_49_), .ZN(n3625) );
  INV_X4 U1376 ( .A(n3627), .ZN(n3432) );
  OAI221_X2 U1377 ( .B1(n4593), .B2(n3628), .C1(n3629), .C2(n4591), .A(n4588), 
        .ZN(n3627) );
  INV_X4 U1378 ( .A(u4_fract_out_pl1_48_), .ZN(n3628) );
  INV_X4 U1380 ( .A(n3630), .ZN(n3430) );
  OAI221_X2 U1381 ( .B1(n4593), .B2(n3631), .C1(n2522), .C2(n4591), .A(n4588), 
        .ZN(n3630) );
  INV_X4 U1382 ( .A(u4_fract_out_pl1_47_), .ZN(n3631) );
  INV_X4 U1384 ( .A(n3632), .ZN(n3431) );
  OAI221_X2 U1385 ( .B1(n4593), .B2(n3633), .C1(n2523), .C2(n4591), .A(n4588), 
        .ZN(n3632) );
  INV_X4 U1386 ( .A(u4_fract_out_pl1_46_), .ZN(n3633) );
  INV_X4 U1388 ( .A(n3419), .ZN(n3614) );
  OAI221_X2 U1389 ( .B1(n4593), .B2(n3634), .C1(n2524), .C2(n4591), .A(n4588), 
        .ZN(n3419) );
  INV_X4 U1390 ( .A(u4_fract_out_pl1_45_), .ZN(n3634) );
  INV_X4 U1392 ( .A(n3421), .ZN(n3601) );
  OAI221_X2 U1393 ( .B1(n4593), .B2(n3635), .C1(n3636), .C2(n4591), .A(n4587), 
        .ZN(n3421) );
  INV_X4 U1394 ( .A(u4_fract_out_pl1_44_), .ZN(n3635) );
  INV_X4 U1396 ( .A(n3420), .ZN(n3600) );
  OAI221_X2 U1397 ( .B1(n4594), .B2(n3637), .C1(n3638), .C2(n4590), .A(n4588), 
        .ZN(n3420) );
  INV_X4 U1398 ( .A(u4_fract_out_pl1_43_), .ZN(n3637) );
  INV_X4 U1400 ( .A(n3639), .ZN(n3422) );
  OAI221_X2 U1401 ( .B1(n4594), .B2(n3640), .C1(n3641), .C2(n4590), .A(n4588), 
        .ZN(n3639) );
  INV_X4 U1402 ( .A(u4_fract_out_pl1_42_), .ZN(n3640) );
  INV_X4 U1404 ( .A(n3642), .ZN(n3423) );
  OAI221_X2 U1405 ( .B1(n4594), .B2(n3643), .C1(n3644), .C2(n4590), .A(n4588), 
        .ZN(n3642) );
  INV_X4 U1406 ( .A(u4_fract_out_pl1_41_), .ZN(n3643) );
  INV_X4 U1408 ( .A(n3645), .ZN(n3424) );
  OAI221_X2 U1409 ( .B1(n4594), .B2(n3646), .C1(n2525), .C2(n4590), .A(n4588), 
        .ZN(n3645) );
  INV_X4 U1410 ( .A(u4_fract_out_pl1_40_), .ZN(n3646) );
  INV_X4 U1412 ( .A(n3647), .ZN(n3425) );
  OAI221_X2 U1413 ( .B1(n4594), .B2(n3648), .C1(n2527), .C2(n4590), .A(n4588), 
        .ZN(n3647) );
  INV_X4 U1414 ( .A(u4_fract_out_pl1_39_), .ZN(n3648) );
  INV_X4 U1416 ( .A(n3412), .ZN(n3602) );
  OAI221_X2 U1417 ( .B1(n4594), .B2(n3649), .C1(n3650), .C2(n4590), .A(n4588), 
        .ZN(n3412) );
  INV_X4 U1418 ( .A(u4_fract_out_pl1_38_), .ZN(n3649) );
  INV_X4 U1420 ( .A(n3414), .ZN(n3603) );
  OAI221_X2 U1421 ( .B1(n4594), .B2(n3651), .C1(n3652), .C2(n4590), .A(n4588), 
        .ZN(n3414) );
  INV_X4 U1422 ( .A(u4_fract_out_pl1_37_), .ZN(n3651) );
  INV_X4 U1424 ( .A(n3413), .ZN(n3604) );
  OAI221_X2 U1425 ( .B1(n4594), .B2(n3653), .C1(n3654), .C2(n4590), .A(n4588), 
        .ZN(n3413) );
  INV_X4 U1426 ( .A(u4_fract_out_pl1_36_), .ZN(n3653) );
  INV_X4 U1428 ( .A(n3655), .ZN(n3417) );
  OAI221_X2 U1429 ( .B1(n4594), .B2(n3656), .C1(n2528), .C2(n4590), .A(n4588), 
        .ZN(n3655) );
  INV_X4 U1430 ( .A(u4_fract_out_pl1_35_), .ZN(n3656) );
  INV_X4 U1432 ( .A(n3657), .ZN(n3415) );
  OAI221_X2 U1433 ( .B1(n4594), .B2(n3658), .C1(n2529), .C2(n4590), .A(n4588), 
        .ZN(n3657) );
  INV_X4 U1434 ( .A(u4_fract_out_pl1_34_), .ZN(n3658) );
  INV_X4 U1436 ( .A(n3659), .ZN(n3416) );
  OAI221_X2 U1437 ( .B1(n4594), .B2(n3660), .C1(n2530), .C2(n4590), .A(n4588), 
        .ZN(n3659) );
  INV_X4 U1438 ( .A(u4_fract_out_pl1_33_), .ZN(n3660) );
  INV_X4 U1440 ( .A(n3404), .ZN(n3605) );
  OAI221_X2 U1441 ( .B1(n4593), .B2(n3661), .C1(n3662), .C2(n4589), .A(n4587), 
        .ZN(n3404) );
  INV_X4 U1442 ( .A(u4_fract_out_pl1_32_), .ZN(n3661) );
  INV_X4 U1444 ( .A(n3406), .ZN(n3606) );
  OAI221_X2 U1445 ( .B1(n4593), .B2(n3663), .C1(n3664), .C2(n4589), .A(n4587), 
        .ZN(n3406) );
  INV_X4 U1446 ( .A(u4_fract_out_pl1_31_), .ZN(n3663) );
  INV_X4 U1448 ( .A(n3405), .ZN(n3607) );
  OAI221_X2 U1449 ( .B1(n4593), .B2(n3665), .C1(n3666), .C2(n4589), .A(n4587), 
        .ZN(n3405) );
  INV_X4 U1450 ( .A(u4_fract_out_pl1_30_), .ZN(n3665) );
  INV_X4 U1452 ( .A(n3667), .ZN(n3407) );
  OAI221_X2 U1453 ( .B1(n4593), .B2(n3668), .C1(n2531), .C2(n4589), .A(n4587), 
        .ZN(n3667) );
  INV_X4 U1454 ( .A(u4_fract_out_pl1_29_), .ZN(n3668) );
  INV_X4 U1456 ( .A(n3669), .ZN(n3408) );
  OAI221_X2 U1457 ( .B1(n4593), .B2(n3670), .C1(n2532), .C2(n4589), .A(n4587), 
        .ZN(n3669) );
  INV_X4 U1458 ( .A(u4_fract_out_pl1_28_), .ZN(n3670) );
  INV_X4 U1460 ( .A(n3671), .ZN(n3409) );
  OAI221_X2 U1461 ( .B1(n4593), .B2(n3672), .C1(n2533), .C2(n4589), .A(n4587), 
        .ZN(n3671) );
  INV_X4 U1462 ( .A(u4_fract_out_pl1_27_), .ZN(n3672) );
  INV_X4 U1464 ( .A(n3673), .ZN(n3410) );
  OAI221_X2 U1465 ( .B1(n4593), .B2(n3674), .C1(n3675), .C2(n4589), .A(n4587), 
        .ZN(n3673) );
  INV_X4 U1466 ( .A(u4_fract_out_pl1_26_), .ZN(n3674) );
  INV_X4 U1468 ( .A(n3448), .ZN(n3590) );
  OAI221_X2 U1469 ( .B1(n4593), .B2(n3676), .C1(n3677), .C2(n4589), .A(n4587), 
        .ZN(n3448) );
  INV_X4 U1470 ( .A(u4_fract_out_pl1_25_), .ZN(n3676) );
  INV_X4 U1472 ( .A(n3450), .ZN(n3591) );
  OAI221_X2 U1473 ( .B1(n4593), .B2(n3678), .C1(n3679), .C2(n4589), .A(n4587), 
        .ZN(n3450) );
  INV_X4 U1474 ( .A(u4_fract_out_pl1_24_), .ZN(n3678) );
  INV_X4 U1476 ( .A(n3449), .ZN(n3592) );
  OAI221_X2 U1477 ( .B1(n4593), .B2(n3680), .C1(n2534), .C2(n4589), .A(n4587), 
        .ZN(n3449) );
  INV_X4 U1478 ( .A(u4_fract_out_pl1_23_), .ZN(n3680) );
  INV_X4 U1480 ( .A(n3681), .ZN(n3453) );
  OAI221_X2 U1481 ( .B1(n4593), .B2(n3682), .C1(n2535), .C2(n4589), .A(n4587), 
        .ZN(n3681) );
  INV_X4 U1482 ( .A(u4_fract_out_pl1_22_), .ZN(n3682) );
  INV_X4 U1484 ( .A(n3683), .ZN(n3451) );
  OAI221_X2 U1485 ( .B1(n4594), .B2(n3684), .C1(n2536), .C2(n4591), .A(n4586), 
        .ZN(n3683) );
  INV_X4 U1486 ( .A(u4_fract_out_pl1_21_), .ZN(n3684) );
  INV_X4 U1488 ( .A(n3685), .ZN(n3452) );
  OAI221_X2 U1489 ( .B1(n4592), .B2(n3686), .C1(n3687), .C2(n4591), .A(n4586), 
        .ZN(n3685) );
  INV_X4 U1490 ( .A(u4_fract_out_pl1_20_), .ZN(n3686) );
  INV_X4 U1492 ( .A(n3440), .ZN(n3593) );
  OAI221_X2 U1493 ( .B1(n4592), .B2(n3688), .C1(n3689), .C2(n4591), .A(n4586), 
        .ZN(n3440) );
  INV_X4 U1494 ( .A(u4_fract_out_pl1_19_), .ZN(n3688) );
  INV_X4 U1496 ( .A(n3442), .ZN(n3594) );
  OAI221_X2 U1497 ( .B1(n4594), .B2(n3690), .C1(n3691), .C2(n4591), .A(n4586), 
        .ZN(n3442) );
  INV_X4 U1498 ( .A(u4_fract_out_pl1_18_), .ZN(n3690) );
  INV_X4 U1500 ( .A(n3441), .ZN(n3595) );
  OAI221_X2 U1501 ( .B1(n4592), .B2(n3692), .C1(n2537), .C2(n4589), .A(n4586), 
        .ZN(n3441) );
  INV_X4 U1502 ( .A(u4_fract_out_pl1_17_), .ZN(n3692) );
  INV_X4 U1504 ( .A(n3693), .ZN(n3443) );
  OAI221_X2 U1505 ( .B1(n4592), .B2(n3694), .C1(n2538), .C2(n4589), .A(n4586), 
        .ZN(n3693) );
  INV_X4 U1506 ( .A(u4_fract_out_pl1_16_), .ZN(n3694) );
  INV_X4 U1508 ( .A(n3695), .ZN(n3444) );
  OAI221_X2 U1509 ( .B1(n4592), .B2(n3696), .C1(n2539), .C2(n4589), .A(n4586), 
        .ZN(n3695) );
  INV_X4 U1510 ( .A(u4_fract_out_pl1_15_), .ZN(n3696) );
  INV_X4 U1512 ( .A(n3697), .ZN(n3445) );
  OAI221_X2 U1513 ( .B1(n4594), .B2(n3698), .C1(n3699), .C2(n4591), .A(n4586), 
        .ZN(n3697) );
  INV_X4 U1514 ( .A(u4_fract_out_pl1_14_), .ZN(n3698) );
  INV_X4 U1516 ( .A(n3700), .ZN(n3446) );
  OAI221_X2 U1517 ( .B1(n4594), .B2(n3701), .C1(n3702), .C2(n4591), .A(n4586), 
        .ZN(n3700) );
  INV_X4 U1518 ( .A(u4_fract_out_pl1_13_), .ZN(n3701) );
  INV_X4 U1520 ( .A(n3334), .ZN(n3578) );
  OAI221_X2 U1521 ( .B1(n4594), .B2(n3703), .C1(n3704), .C2(n4591), .A(n4586), 
        .ZN(n3334) );
  INV_X4 U1522 ( .A(u4_fract_out_pl1_12_), .ZN(n3703) );
  INV_X4 U1524 ( .A(n3336), .ZN(n3579) );
  OAI221_X2 U1525 ( .B1(n4594), .B2(n3705), .C1(n2540), .C2(n4591), .A(n4586), 
        .ZN(n3336) );
  INV_X4 U1526 ( .A(u4_fract_out_pl1_11_), .ZN(n3705) );
  INV_X4 U1528 ( .A(n3335), .ZN(n3580) );
  OAI221_X2 U1529 ( .B1(n4592), .B2(n3706), .C1(n2541), .C2(n4590), .A(n4586), 
        .ZN(n3335) );
  INV_X4 U1530 ( .A(u4_fract_out_pl1_10_), .ZN(n3706) );
  INV_X4 U1532 ( .A(n3707), .ZN(n3337) );
  OAI221_X2 U1533 ( .B1(n4592), .B2(n3708), .C1(n3709), .C2(n4591), .A(n4586), 
        .ZN(n3707) );
  INV_X4 U1534 ( .A(u4_fract_out_pl1_9_), .ZN(n3708) );
  INV_X4 U1536 ( .A(n3710), .ZN(n3338) );
  OAI221_X2 U1537 ( .B1(n4592), .B2(n3711), .C1(n3712), .C2(n4589), .A(n4586), 
        .ZN(n3710) );
  INV_X4 U1538 ( .A(u4_fract_out_pl1_8_), .ZN(n3711) );
  INV_X4 U1540 ( .A(n3713), .ZN(n3339) );
  OAI221_X2 U1541 ( .B1(n4592), .B2(n3714), .C1(n3715), .C2(n4591), .A(n4586), 
        .ZN(n3713) );
  INV_X4 U1542 ( .A(u4_fract_out_pl1_7_), .ZN(n3714) );
  INV_X4 U1544 ( .A(n3436), .ZN(n3340) );
  OAI221_X2 U1545 ( .B1(n4592), .B2(n3716), .C1(n3717), .C2(n4590), .A(n4586), 
        .ZN(n3436) );
  INV_X4 U1546 ( .A(u4_fract_out_pl1_6_), .ZN(n3716) );
  INV_X4 U1548 ( .A(n3326), .ZN(n3581) );
  OAI221_X2 U1549 ( .B1(n4592), .B2(n3718), .C1(n2519), .C2(n4590), .A(n4586), 
        .ZN(n3326) );
  INV_X4 U1550 ( .A(u4_fract_out_pl1_5_), .ZN(n3718) );
  INV_X4 U1552 ( .A(n3328), .ZN(n3582) );
  OAI221_X2 U1553 ( .B1(n4592), .B2(n3719), .C1(n3720), .C2(n4590), .A(n4586), 
        .ZN(n3328) );
  INV_X4 U1554 ( .A(u4_fract_out_pl1_4_), .ZN(n3719) );
  INV_X4 U1556 ( .A(n3327), .ZN(n3437) );
  OAI221_X2 U1557 ( .B1(n4592), .B2(n3721), .C1(n2526), .C2(n4590), .A(n4586), 
        .ZN(n3327) );
  INV_X4 U1558 ( .A(u4_fract_out_pl1_3_), .ZN(n3721) );
  INV_X4 U1560 ( .A(n3722), .ZN(n3329) );
  OAI221_X2 U1561 ( .B1(n4592), .B2(n3723), .C1(n3724), .C2(n4589), .A(n4586), 
        .ZN(n3722) );
  INV_X4 U1562 ( .A(u4_fract_out_pl1_2_), .ZN(n3723) );
  INV_X4 U1564 ( .A(n3725), .ZN(n3330) );
  OAI221_X2 U1565 ( .B1(n4592), .B2(n3726), .C1(n3727), .C2(n4590), .A(n4586), 
        .ZN(n3725) );
  INV_X4 U1566 ( .A(u4_fract_out_pl1_1_), .ZN(n3726) );
  OAI22_X2 U1567 ( .A1(n6310), .A2(n3331), .B1(n3341), .B2(n3619), .ZN(N793)
         );
  OAI22_X2 U1569 ( .A1(n3308), .A2(n4355), .B1(n2507), .B2(n3468), .ZN(n3728)
         );
  AOI22_X2 U1570 ( .A1(opb_00), .A2(opa_inf), .B1(opb_inf), .B2(opa_00), .ZN(
        n3468) );
  NAND2_X2 U1571 ( .A1(opa_00), .A2(opb_00), .ZN(n3308) );
  INV_X4 U1572 ( .A(n3729), .ZN(n3331) );
  OAI221_X2 U1573 ( .B1(n4592), .B2(n3730), .C1(n3731), .C2(n4590), .A(n4586), 
        .ZN(n3729) );
  OAI221_X2 U1580 ( .B1(n4351), .B2(n3739), .C1(u4_N6410), .C2(n3740), .A(
        n3741), .ZN(n3738) );
  INV_X4 U1581 ( .A(u4_fract_out_pl1_0_), .ZN(n3730) );
  OAI22_X2 U1583 ( .A1(u4_N6410), .A2(n3743), .B1(n3744), .B2(n4351), .ZN(
        n3742) );
  INV_X4 U1584 ( .A(n3739), .ZN(n3744) );
  AND3_X2 U1585 ( .A1(n3745), .A2(n3552), .A3(n3554), .ZN(n3734) );
  AND4_X2 U1587 ( .A1(n3584), .A2(n3583), .A3(n3746), .A4(n3747), .ZN(n3332)
         );
  NOR4_X2 U1588 ( .A1(n3748), .A2(n3389), .A3(n3617), .A4(n3388), .ZN(n3747)
         );
  INV_X4 U1593 ( .A(n3615), .ZN(n3393) );
  INV_X4 U1595 ( .A(n3539), .ZN(n3395) );
  INV_X4 U1597 ( .A(n3540), .ZN(n3394) );
  INV_X4 U1600 ( .A(n3534), .ZN(n3398) );
  INV_X4 U1604 ( .A(n3585), .ZN(n3618) );
  NAND2_X2 U1608 ( .A1(n6315), .A2(n3765), .ZN(n3758) );
  NAND2_X2 U1609 ( .A1(n3761), .A2(n6315), .ZN(n3757) );
  NAND2_X2 U1610 ( .A1(n3745), .A2(n3766), .ZN(n3760) );
  OAI211_X2 U1614 ( .C1(n3769), .C2(n3556), .A(u4_N6410), .B(n3297), .ZN(n3768) );
  AND4_X2 U1615 ( .A1(n3770), .A2(n6466), .A3(u4_N6249), .A4(n3771), .ZN(n3769) );
  OR4_X2 U1616 ( .A1(u4_exp_out_0_), .A2(u4_exp_out_8_), .A3(u4_exp_out_9_), 
        .A4(n3772), .ZN(n3770) );
  AND4_X2 U1618 ( .A1(sign), .A2(rmode_r3[1]), .A3(n3775), .A4(n4452), .ZN(
        n3774) );
  OAI221_X2 U1619 ( .B1(n3776), .B2(n2514), .C1(n3777), .C2(n4653), .A(n3778), 
        .ZN(n3775) );
  NAND4_X2 U1620 ( .A1(n3762), .A2(n4656), .A3(n3779), .A4(n3780), .ZN(n3778)
         );
  OR4_X2 U1621 ( .A1(n3772), .A2(n2450), .A3(n2443), .A4(u4_exp_out_mi1[0]), 
        .ZN(n3779) );
  INV_X4 U1623 ( .A(u4_exp_out_9_), .ZN(n2443) );
  NAND2_X2 U1624 ( .A1(n3781), .A2(n3782), .ZN(n3772) );
  NOR4_X2 U1625 ( .A1(u4_exp_out_10_), .A2(n2453), .A3(n2456), .A4(n2459), 
        .ZN(n3782) );
  NOR4_X2 U1626 ( .A1(n2462), .A2(n2465), .A3(n2468), .A4(n2471), .ZN(n3781)
         );
  OAI211_X2 U1630 ( .C1(n4355), .C2(n3481), .A(n6306), .B(n3554), .ZN(n3765)
         );
  INV_X4 U1631 ( .A(n3478), .ZN(n3554) );
  AOI22_X2 U1632 ( .A1(n4540), .A2(n3785), .B1(n3786), .B2(n3297), .ZN(n3784)
         );
  NAND4_X2 U1636 ( .A1(u4_N6249), .A2(n6466), .A3(n3791), .A4(n3488), .ZN(
        n3790) );
  NAND4_X2 U1637 ( .A1(n3762), .A2(n3763), .A3(n3792), .A4(n3793), .ZN(n3791)
         );
  AND4_X2 U1638 ( .A1(n3794), .A2(n3752), .A3(n3751), .A4(n3749), .ZN(n3793)
         );
  OAI211_X2 U1639 ( .C1(n3795), .C2(n2465), .A(n3796), .B(n3797), .ZN(n3749)
         );
  AOI221_X2 U1640 ( .B1(u4_exp_fix_divb[3]), .B2(n3798), .C1(
        u4_exp_fix_diva[3]), .C2(n3799), .A(n3800), .ZN(n3797) );
  INV_X4 U1641 ( .A(n3801), .ZN(n3800) );
  AOI22_X2 U1642 ( .A1(u4_exp_next_mi_3_), .A2(n3802), .B1(exp_r[3]), .B2(
        n3803), .ZN(n3801) );
  AOI22_X2 U1643 ( .A1(u4_exp_out_mi1[3]), .A2(n3804), .B1(u4_exp_out_pl1_3_), 
        .B2(n3805), .ZN(n3796) );
  OAI211_X2 U1644 ( .C1(n3795), .C2(n2462), .A(n3806), .B(n3807), .ZN(n3751)
         );
  AOI221_X2 U1645 ( .B1(u4_exp_fix_divb[4]), .B2(n3798), .C1(
        u4_exp_fix_diva[4]), .C2(n3799), .A(n3808), .ZN(n3807) );
  INV_X4 U1646 ( .A(n3809), .ZN(n3808) );
  AOI22_X2 U1647 ( .A1(u4_exp_next_mi_4_), .A2(n3802), .B1(n4282), .B2(n3803), 
        .ZN(n3809) );
  AOI22_X2 U1648 ( .A1(u4_exp_out_mi1[4]), .A2(n3804), .B1(u4_exp_out_pl1_4_), 
        .B2(n3805), .ZN(n3806) );
  OAI211_X2 U1649 ( .C1(n3795), .C2(n2468), .A(n3810), .B(n3811), .ZN(n3752)
         );
  AOI221_X2 U1650 ( .B1(u4_exp_fix_divb[2]), .B2(n3798), .C1(
        u4_exp_fix_diva[2]), .C2(n3799), .A(n3812), .ZN(n3811) );
  INV_X4 U1651 ( .A(n3813), .ZN(n3812) );
  AOI22_X2 U1652 ( .A1(u4_exp_next_mi_2_), .A2(n3802), .B1(n4315), .B2(n3803), 
        .ZN(n3813) );
  AOI22_X2 U1653 ( .A1(u4_exp_out_mi1[2]), .A2(n3804), .B1(u4_exp_out_pl1_2_), 
        .B2(n3805), .ZN(n3810) );
  INV_X4 U1654 ( .A(u4_exp_out_2_), .ZN(n2468) );
  AND3_X2 U1655 ( .A1(n3755), .A2(n3754), .A3(n3753), .ZN(n3794) );
  OAI211_X2 U1656 ( .C1(n3795), .C2(n2459), .A(n3814), .B(n3815), .ZN(n3753)
         );
  AOI221_X2 U1657 ( .B1(u4_exp_fix_divb[5]), .B2(n3798), .C1(
        u4_exp_fix_diva[5]), .C2(n3799), .A(n3816), .ZN(n3815) );
  INV_X4 U1658 ( .A(n3817), .ZN(n3816) );
  AOI22_X2 U1659 ( .A1(u4_exp_next_mi_5_), .A2(n3802), .B1(n4290), .B2(n3803), 
        .ZN(n3817) );
  AOI22_X2 U1660 ( .A1(u4_exp_out_mi1[5]), .A2(n3804), .B1(u4_exp_out_pl1_5_), 
        .B2(n3805), .ZN(n3814) );
  OAI211_X2 U1661 ( .C1(n3795), .C2(n2453), .A(n3818), .B(n3819), .ZN(n3754)
         );
  AOI221_X2 U1662 ( .B1(u4_exp_fix_divb[7]), .B2(n3798), .C1(
        u4_exp_fix_diva[7]), .C2(n3799), .A(n3820), .ZN(n3819) );
  INV_X4 U1663 ( .A(n3821), .ZN(n3820) );
  AOI22_X2 U1664 ( .A1(u4_exp_next_mi_7_), .A2(n3802), .B1(n4281), .B2(n3803), 
        .ZN(n3821) );
  AOI22_X2 U1665 ( .A1(u4_exp_out_mi1[7]), .A2(n3804), .B1(u4_exp_out_pl1_7_), 
        .B2(n3805), .ZN(n3818) );
  OAI211_X2 U1666 ( .C1(n3795), .C2(n2456), .A(n3822), .B(n3823), .ZN(n3755)
         );
  AOI221_X2 U1667 ( .B1(u4_exp_fix_divb[6]), .B2(n3798), .C1(
        u4_exp_fix_diva[6]), .C2(n3799), .A(n3824), .ZN(n3823) );
  INV_X4 U1668 ( .A(n3825), .ZN(n3824) );
  AOI22_X2 U1669 ( .A1(u4_exp_next_mi_6_), .A2(n3802), .B1(exp_r[6]), .B2(
        n3803), .ZN(n3825) );
  AOI22_X2 U1670 ( .A1(u4_exp_out_mi1[6]), .A2(n3804), .B1(u4_exp_out_pl1_6_), 
        .B2(n3805), .ZN(n3822) );
  AND3_X2 U1671 ( .A1(n3764), .A2(n3759), .A3(n3756), .ZN(n3792) );
  AND3_X2 U1672 ( .A1(n3826), .A2(n3827), .A3(n3828), .ZN(n3756) );
  AOI22_X2 U1674 ( .A1(u4_exp_fix_divb[0]), .A2(n3798), .B1(u4_exp_fix_diva[0]), .B2(n3799), .ZN(n3827) );
  AOI22_X2 U1675 ( .A1(u4_exp_out_mi1[0]), .A2(n3804), .B1(n3803), .B2(n4600), 
        .ZN(n3826) );
  OAI211_X2 U1676 ( .C1(n3795), .C2(n2471), .A(n3830), .B(n3831), .ZN(n3759)
         );
  AOI221_X2 U1677 ( .B1(u4_exp_fix_divb[1]), .B2(n3798), .C1(
        u4_exp_fix_diva[1]), .C2(n3799), .A(n3832), .ZN(n3831) );
  INV_X4 U1678 ( .A(n3833), .ZN(n3832) );
  AOI22_X2 U1679 ( .A1(u4_exp_next_mi_1_), .A2(n3802), .B1(exp_r[1]), .B2(
        n3803), .ZN(n3833) );
  AOI22_X2 U1680 ( .A1(u4_exp_out_mi1[1]), .A2(n3804), .B1(u4_exp_out_pl1_1_), 
        .B2(n3805), .ZN(n3830) );
  INV_X4 U1681 ( .A(u4_exp_out_1_), .ZN(n2471) );
  INV_X4 U1683 ( .A(n3836), .ZN(n3835) );
  AND3_X2 U1684 ( .A1(n3837), .A2(n3838), .A3(n3839), .ZN(n3763) );
  AOI22_X2 U1686 ( .A1(u4_exp_fix_divb[9]), .A2(n3798), .B1(u4_exp_fix_diva[9]), .B2(n3799), .ZN(n3838) );
  AOI22_X2 U1687 ( .A1(u4_exp_out_mi1[9]), .A2(n3804), .B1(n3803), .B2(n4289), 
        .ZN(n3837) );
  AND3_X2 U1688 ( .A1(n3840), .A2(n3841), .A3(n3842), .ZN(n3762) );
  AOI22_X2 U1690 ( .A1(u4_exp_fix_divb[10]), .A2(n3798), .B1(
        u4_exp_fix_diva[10]), .B2(n3799), .ZN(n3841) );
  AOI22_X2 U1691 ( .A1(u4_exp_out_mi1[10]), .A2(n3804), .B1(n3803), .B2(n4656), 
        .ZN(n3840) );
  OAI22_X2 U1695 ( .A1(opas_r2), .A2(n6467), .B1(n6308), .B2(n3843), .ZN(n2435) );
  NAND2_X2 U1696 ( .A1(n3556), .A2(n4823), .ZN(n3481) );
  AND3_X2 U1698 ( .A1(n3844), .A2(n3845), .A3(n3846), .ZN(n3764) );
  INV_X4 U1701 ( .A(n3848), .ZN(n2440) );
  NAND2_X2 U1703 ( .A1(n3836), .A2(n3850), .ZN(n3829) );
  AOI22_X2 U1706 ( .A1(n4823), .A2(n3847), .B1(n6305), .B2(n3852), .ZN(n3836)
         );
  INV_X4 U1708 ( .A(n3551), .ZN(n3557) );
  NAND2_X2 U1709 ( .A1(n3740), .A2(u4_fract_out_pl1_52_), .ZN(n3847) );
  INV_X4 U1710 ( .A(n3743), .ZN(n3740) );
  AOI22_X2 U1712 ( .A1(u4_exp_fix_divb[8]), .A2(n3798), .B1(u4_exp_fix_diva[8]), .B2(n3799), .ZN(n3845) );
  AOI22_X2 U1716 ( .A1(u4_exp_out_mi1[8]), .A2(n3804), .B1(n3803), .B2(n4353), 
        .ZN(n3844) );
  NAND4_X2 U1718 ( .A1(u4_exp_out_1_), .A2(u4_exp_out_2_), .A3(n3856), .A4(
        n3857), .ZN(n3551) );
  NOR4_X2 U1719 ( .A1(n3858), .A2(n2456), .A3(n2450), .A4(n2453), .ZN(n3857)
         );
  INV_X4 U1720 ( .A(u4_exp_out_7_), .ZN(n2453) );
  INV_X4 U1721 ( .A(u4_exp_out_8_), .ZN(n2450) );
  INV_X4 U1722 ( .A(u4_exp_out_6_), .ZN(n2456) );
  INV_X4 U1725 ( .A(u4_exp_out_4_), .ZN(n2462) );
  INV_X4 U1726 ( .A(u4_exp_out_5_), .ZN(n2459) );
  INV_X4 U1727 ( .A(u4_exp_out_3_), .ZN(n2465) );
  AND4_X2 U1728 ( .A1(n3854), .A2(n6466), .A3(u4_fract_out_0_), .A4(n3853), 
        .ZN(n3849) );
  INV_X4 U1729 ( .A(n3731), .ZN(u4_fract_out_0_) );
  NAND4_X2 U1730 ( .A1(n4289), .A2(n4600), .A3(n3859), .A4(n3860), .ZN(n3787)
         );
  NOR4_X2 U1731 ( .A1(n3861), .A2(n4299), .A3(n4317), .A4(n4347), .ZN(n3860)
         );
  AND3_X2 U1733 ( .A1(exp_r[1]), .A2(n4655), .A3(n4315), .ZN(n3859) );
  NAND2_X2 U1736 ( .A1(u4_fract_out_pl1_52_), .A2(n3739), .ZN(n3834) );
  OAI211_X2 U1738 ( .C1(n3864), .C2(n3485), .A(n4441), .B(n6342), .ZN(n3863)
         );
  NAND2_X2 U1739 ( .A1(n3865), .A2(n3866), .ZN(n3485) );
  NAND4_X2 U1744 ( .A1(n6404), .A2(n6403), .A3(n2763), .A4(n3872), .ZN(n3869)
         );
  NOR4_X2 U1746 ( .A1(n3874), .A2(n3875), .A3(n2634), .A4(n2771), .ZN(n3867)
         );
  OR3_X2 U1747 ( .A1(n2635), .A2(n2561), .A3(n2604), .ZN(n3875) );
  NAND4_X2 U1748 ( .A1(n3876), .A2(n2636), .A3(n3877), .A4(n3878), .ZN(n3874)
         );
  AND4_X2 U1751 ( .A1(u4_N6917), .A2(n6317), .A3(n3544), .A4(n2434), .ZN(n3881) );
  OAI211_X2 U1754 ( .C1(n4540), .C2(n3488), .A(n3473), .B(n3882), .ZN(n3885)
         );
  NAND2_X2 U1755 ( .A1(n3886), .A2(n3887), .ZN(n3473) );
  NOR4_X2 U1756 ( .A1(n3888), .A2(n3889), .A3(n3890), .A4(n3891), .ZN(n3887)
         );
  NAND4_X2 U1757 ( .A1(n2529), .A2(n2528), .A3(n2530), .A4(n3892), .ZN(n3891)
         );
  INV_X4 U1759 ( .A(n3652), .ZN(u4_fract_out_37_) );
  AOI22_X2 U1760 ( .A1(u4_N5997), .A2(n4578), .B1(u4_N6105), .B2(n4576), .ZN(
        n3652) );
  INV_X4 U1761 ( .A(n3650), .ZN(u4_fract_out_38_) );
  AOI22_X2 U1762 ( .A1(u4_N5998), .A2(n4582), .B1(u4_N6106), .B2(n4577), .ZN(
        n3650) );
  INV_X4 U1763 ( .A(n3654), .ZN(u4_fract_out_36_) );
  AOI22_X2 U1764 ( .A1(u4_N5996), .A2(n4582), .B1(u4_N6104), .B2(n4577), .ZN(
        n3654) );
  AOI22_X2 U1765 ( .A1(u4_N5993), .A2(n4582), .B1(u4_N6101), .B2(n4577), .ZN(
        n2530) );
  AOI22_X2 U1766 ( .A1(u4_N5995), .A2(n4582), .B1(u4_N6103), .B2(n4577), .ZN(
        n2528) );
  AOI22_X2 U1767 ( .A1(u4_N5994), .A2(n4582), .B1(u4_N6102), .B2(n4577), .ZN(
        n2529) );
  NAND4_X2 U1768 ( .A1(n2526), .A2(n2525), .A3(n2527), .A4(n3895), .ZN(n3890)
         );
  NOR4_X2 U1769 ( .A1(u4_fract_out_44_), .A2(u4_fract_out_43_), .A3(
        u4_fract_out_42_), .A4(u4_fract_out_41_), .ZN(n3895) );
  INV_X4 U1770 ( .A(n3644), .ZN(u4_fract_out_41_) );
  AOI22_X2 U1771 ( .A1(u4_N6001), .A2(n4582), .B1(u4_N6109), .B2(n4577), .ZN(
        n3644) );
  INV_X4 U1772 ( .A(n3641), .ZN(u4_fract_out_42_) );
  AOI22_X2 U1773 ( .A1(u4_N6002), .A2(n4582), .B1(u4_N6110), .B2(n4577), .ZN(
        n3641) );
  INV_X4 U1774 ( .A(n3638), .ZN(u4_fract_out_43_) );
  AOI22_X2 U1775 ( .A1(u4_N6003), .A2(n4582), .B1(u4_N6111), .B2(n4577), .ZN(
        n3638) );
  INV_X4 U1776 ( .A(n3636), .ZN(u4_fract_out_44_) );
  AOI22_X2 U1777 ( .A1(u4_N6004), .A2(n4582), .B1(u4_N6112), .B2(n4577), .ZN(
        n3636) );
  AOI22_X2 U1778 ( .A1(u4_N5999), .A2(n4582), .B1(u4_N6107), .B2(n4577), .ZN(
        n2527) );
  AOI22_X2 U1779 ( .A1(u4_N6000), .A2(n4581), .B1(u4_N6108), .B2(n4577), .ZN(
        n2525) );
  AOI22_X2 U1780 ( .A1(u4_N5963), .A2(n4581), .B1(u4_N6071), .B2(n4577), .ZN(
        n2526) );
  NAND4_X2 U1781 ( .A1(n2523), .A2(n2522), .A3(n2524), .A4(n3896), .ZN(n3889)
         );
  INV_X4 U1783 ( .A(n3626), .ZN(u4_fract_out_49_) );
  AOI22_X2 U1784 ( .A1(u4_N6009), .A2(n4581), .B1(u4_N6117), .B2(n4577), .ZN(
        n3626) );
  INV_X4 U1785 ( .A(n3720), .ZN(u4_fract_out_4_) );
  AOI22_X2 U1786 ( .A1(u4_N5964), .A2(n4581), .B1(u4_N6072), .B2(n4577), .ZN(
        n3720) );
  INV_X4 U1787 ( .A(n3629), .ZN(u4_fract_out_48_) );
  AOI22_X2 U1788 ( .A1(u4_N6008), .A2(n4581), .B1(u4_N6116), .B2(n4577), .ZN(
        n3629) );
  AOI22_X2 U1789 ( .A1(u4_N6005), .A2(n4581), .B1(u4_N6113), .B2(n4577), .ZN(
        n2524) );
  AOI22_X2 U1790 ( .A1(u4_N6007), .A2(n4581), .B1(u4_N6115), .B2(n4577), .ZN(
        n2522) );
  AOI22_X2 U1791 ( .A1(u4_N6006), .A2(n4581), .B1(u4_N6114), .B2(n4577), .ZN(
        n2523) );
  NAND4_X2 U1792 ( .A1(n2520), .A2(n2519), .A3(n2521), .A4(n3897), .ZN(n3888)
         );
  NOR4_X2 U1793 ( .A1(u4_fract_out_9_), .A2(u4_fract_out_8_), .A3(
        u4_fract_out_7_), .A4(u4_fract_out_6_), .ZN(n3897) );
  INV_X4 U1794 ( .A(n3717), .ZN(u4_fract_out_6_) );
  AOI22_X2 U1795 ( .A1(u4_N5966), .A2(n4581), .B1(u4_N6074), .B2(n4577), .ZN(
        n3717) );
  INV_X4 U1796 ( .A(n3715), .ZN(u4_fract_out_7_) );
  AOI22_X2 U1797 ( .A1(u4_N5967), .A2(n4581), .B1(u4_N6075), .B2(n4577), .ZN(
        n3715) );
  INV_X4 U1798 ( .A(n3712), .ZN(u4_fract_out_8_) );
  AOI22_X2 U1799 ( .A1(u4_N5968), .A2(n4581), .B1(u4_N6076), .B2(n3894), .ZN(
        n3712) );
  INV_X4 U1800 ( .A(n3709), .ZN(u4_fract_out_9_) );
  AOI22_X2 U1801 ( .A1(u4_N5969), .A2(n4580), .B1(u4_N6077), .B2(n3894), .ZN(
        n3709) );
  AOI22_X2 U1802 ( .A1(u4_N6010), .A2(n4580), .B1(u4_N6118), .B2(n3894), .ZN(
        n2521) );
  AOI22_X2 U1803 ( .A1(u4_N5965), .A2(n4580), .B1(u4_N6073), .B2(n3894), .ZN(
        n2519) );
  AOI22_X2 U1804 ( .A1(u4_N6011), .A2(n4580), .B1(u4_N6119), .B2(n3894), .ZN(
        n2520) );
  NOR4_X2 U1805 ( .A1(n3898), .A2(n3899), .A3(n3900), .A4(n3901), .ZN(n3886)
         );
  NAND4_X2 U1806 ( .A1(n2541), .A2(n2540), .A3(n3731), .A4(n3902), .ZN(n3901)
         );
  INV_X4 U1808 ( .A(n3702), .ZN(u4_fract_out_13_) );
  AOI22_X2 U1809 ( .A1(u4_N5973), .A2(n4580), .B1(u4_N6081), .B2(n3894), .ZN(
        n3702) );
  INV_X4 U1810 ( .A(n3699), .ZN(u4_fract_out_14_) );
  AOI22_X2 U1811 ( .A1(u4_N5974), .A2(n4580), .B1(u4_N6082), .B2(n3894), .ZN(
        n3699) );
  INV_X4 U1812 ( .A(n3704), .ZN(u4_fract_out_12_) );
  AOI22_X2 U1813 ( .A1(u4_N5972), .A2(n4580), .B1(u4_N6080), .B2(n3894), .ZN(
        n3704) );
  AOI22_X2 U1814 ( .A1(u4_N5960), .A2(n4580), .B1(u4_N6068), .B2(n3894), .ZN(
        n3731) );
  AOI22_X2 U1815 ( .A1(u4_N5971), .A2(n4580), .B1(u4_N6079), .B2(n3894), .ZN(
        n2540) );
  AOI22_X2 U1816 ( .A1(u4_N5970), .A2(n4580), .B1(u4_N6078), .B2(n4576), .ZN(
        n2541) );
  NAND4_X2 U1817 ( .A1(n2538), .A2(n2537), .A3(n2539), .A4(n3903), .ZN(n3900)
         );
  NOR4_X2 U1818 ( .A1(u4_fract_out_20_), .A2(u4_fract_out_1_), .A3(
        u4_fract_out_19_), .A4(u4_fract_out_18_), .ZN(n3903) );
  INV_X4 U1819 ( .A(n3691), .ZN(u4_fract_out_18_) );
  AOI22_X2 U1820 ( .A1(u4_N5978), .A2(n4579), .B1(u4_N6086), .B2(n4576), .ZN(
        n3691) );
  INV_X4 U1821 ( .A(n3689), .ZN(u4_fract_out_19_) );
  AOI22_X2 U1822 ( .A1(u4_N5979), .A2(n4579), .B1(u4_N6087), .B2(n4576), .ZN(
        n3689) );
  INV_X4 U1823 ( .A(n3727), .ZN(u4_fract_out_1_) );
  AOI22_X2 U1824 ( .A1(u4_N5961), .A2(n4579), .B1(u4_N6069), .B2(n4576), .ZN(
        n3727) );
  INV_X4 U1825 ( .A(n3687), .ZN(u4_fract_out_20_) );
  AOI22_X2 U1826 ( .A1(u4_N5980), .A2(n4579), .B1(u4_N6088), .B2(n4576), .ZN(
        n3687) );
  AOI22_X2 U1827 ( .A1(u4_N5975), .A2(n4579), .B1(u4_N6083), .B2(n4576), .ZN(
        n2539) );
  AOI22_X2 U1828 ( .A1(u4_N5977), .A2(n4579), .B1(u4_N6085), .B2(n4576), .ZN(
        n2537) );
  AOI22_X2 U1829 ( .A1(u4_N5976), .A2(n4579), .B1(u4_N6084), .B2(n4576), .ZN(
        n2538) );
  NAND4_X2 U1830 ( .A1(n2535), .A2(n2534), .A3(n2536), .A4(n3904), .ZN(n3899)
         );
  INV_X4 U1832 ( .A(n3677), .ZN(u4_fract_out_25_) );
  AOI22_X2 U1833 ( .A1(u4_N5985), .A2(n4579), .B1(u4_N6093), .B2(n4576), .ZN(
        n3677) );
  INV_X4 U1834 ( .A(n3675), .ZN(u4_fract_out_26_) );
  AOI22_X2 U1835 ( .A1(u4_N5986), .A2(n4579), .B1(u4_N6094), .B2(n4576), .ZN(
        n3675) );
  INV_X4 U1836 ( .A(n3679), .ZN(u4_fract_out_24_) );
  AOI22_X2 U1837 ( .A1(u4_N5984), .A2(n4579), .B1(u4_N6092), .B2(n4576), .ZN(
        n3679) );
  AOI22_X2 U1838 ( .A1(u4_N5981), .A2(n4579), .B1(u4_N6089), .B2(n4577), .ZN(
        n2536) );
  AOI22_X2 U1839 ( .A1(u4_N5983), .A2(n4578), .B1(u4_N6091), .B2(n4576), .ZN(
        n2534) );
  AOI22_X2 U1840 ( .A1(u4_N5982), .A2(n4578), .B1(u4_N6090), .B2(n4576), .ZN(
        n2535) );
  NAND4_X2 U1841 ( .A1(n2532), .A2(n2531), .A3(n2533), .A4(n3905), .ZN(n3898)
         );
  NOR4_X2 U1842 ( .A1(u4_fract_out_32_), .A2(u4_fract_out_31_), .A3(
        u4_fract_out_30_), .A4(u4_fract_out_2_), .ZN(n3905) );
  INV_X4 U1843 ( .A(n3724), .ZN(u4_fract_out_2_) );
  AOI22_X2 U1844 ( .A1(u4_N5962), .A2(n4578), .B1(u4_N6070), .B2(n4576), .ZN(
        n3724) );
  INV_X4 U1845 ( .A(n3666), .ZN(u4_fract_out_30_) );
  AOI22_X2 U1846 ( .A1(u4_N5990), .A2(n4578), .B1(u4_N6098), .B2(n4576), .ZN(
        n3666) );
  INV_X4 U1847 ( .A(n3664), .ZN(u4_fract_out_31_) );
  AOI22_X2 U1848 ( .A1(u4_N5991), .A2(n4578), .B1(u4_N6099), .B2(n4577), .ZN(
        n3664) );
  INV_X4 U1849 ( .A(n3662), .ZN(u4_fract_out_32_) );
  AOI22_X2 U1850 ( .A1(u4_N5992), .A2(n4578), .B1(u4_N6100), .B2(n4576), .ZN(
        n3662) );
  AOI22_X2 U1851 ( .A1(u4_N5987), .A2(n4578), .B1(u4_N6095), .B2(n4576), .ZN(
        n2533) );
  AOI22_X2 U1852 ( .A1(u4_N5989), .A2(n4578), .B1(u4_N6097), .B2(n4576), .ZN(
        n2531) );
  AOI22_X2 U1853 ( .A1(u4_N5988), .A2(n4578), .B1(u4_N6096), .B2(n4576), .ZN(
        n2532) );
  OAI22_X2 U1856 ( .A1(exp_ovf_r[0]), .A2(n6095), .B1(exp_ovf_r[1]), .B2(n3780), .ZN(n3906) );
  NAND4_X2 U1857 ( .A1(n4656), .A2(n4349), .A3(n3907), .A4(n3908), .ZN(n3780)
         );
  NOR4_X2 U1858 ( .A1(n3909), .A2(n4282), .A3(exp_r[6]), .A4(n4290), .ZN(n3908) );
  OR3_X2 U1859 ( .A1(n4353), .A2(n4289), .A3(n4281), .ZN(n3909) );
  OR2_X2 U1862 ( .A1(n3853), .A2(n3854), .ZN(n3544) );
  AND4_X2 U1864 ( .A1(u4_N5843), .A2(n6369), .A3(n6352), .A4(n2761), .ZN(n3911) );
  AND4_X2 U1865 ( .A1(n6365), .A2(n6360), .A3(n6359), .A4(n2449), .ZN(n3910)
         );
  AOI22_X2 U1868 ( .A1(n3914), .A2(n4577), .B1(n3915), .B2(n4578), .ZN(n3866)
         );
  OR4_X2 U1869 ( .A1(n3916), .A2(n3917), .A3(n3918), .A4(n3919), .ZN(n3915) );
  NAND4_X2 U1870 ( .A1(n3920), .A2(n3921), .A3(n3922), .A4(n3923), .ZN(n3919)
         );
  NOR4_X2 U1871 ( .A1(u4_N5918), .A2(u4_N5917), .A3(u4_N5916), .A4(u4_N5915), 
        .ZN(n3923) );
  NAND4_X2 U1875 ( .A1(n3924), .A2(n3925), .A3(n3926), .A4(n3927), .ZN(n3918)
         );
  NOR4_X2 U1876 ( .A1(u4_N5931), .A2(u4_N5930), .A3(u4_N5929), .A4(u4_N5928), 
        .ZN(n3927) );
  NAND4_X2 U1880 ( .A1(n3928), .A2(n3929), .A3(n3930), .A4(n3931), .ZN(n3917)
         );
  NOR4_X2 U1881 ( .A1(u4_N5944), .A2(u4_N5943), .A3(u4_N5942), .A4(u4_N5941), 
        .ZN(n3931) );
  NAND4_X2 U1885 ( .A1(n3932), .A2(n3933), .A3(n3934), .A4(n3935), .ZN(n3916)
         );
  NOR4_X2 U1886 ( .A1(u4_N5958), .A2(u4_N5957), .A3(u4_N5956), .A4(u4_N5955), 
        .ZN(n3935) );
  NOR4_X2 U1888 ( .A1(u4_N5951), .A2(u4_N5950), .A3(u4_N5949), .A4(u4_N5948), 
        .ZN(n3933) );
  OR4_X2 U1890 ( .A1(n3936), .A2(n3937), .A3(n3938), .A4(n3939), .ZN(n3914) );
  NAND4_X2 U1891 ( .A1(n3940), .A2(n3941), .A3(n3942), .A4(n3943), .ZN(n3939)
         );
  NOR4_X2 U1892 ( .A1(u4_N6026), .A2(u4_N6025), .A3(u4_N6024), .A4(u4_N6023), 
        .ZN(n3943) );
  NAND4_X2 U1896 ( .A1(n3944), .A2(n3945), .A3(n3946), .A4(n3947), .ZN(n3938)
         );
  NOR4_X2 U1897 ( .A1(u4_N6039), .A2(u4_N6038), .A3(u4_N6037), .A4(u4_N6036), 
        .ZN(n3947) );
  NAND4_X2 U1901 ( .A1(n3948), .A2(n3949), .A3(n3950), .A4(n3951), .ZN(n3937)
         );
  NOR4_X2 U1902 ( .A1(u4_N6052), .A2(u4_N6051), .A3(u4_N6050), .A4(u4_N6049), 
        .ZN(n3951) );
  NAND4_X2 U1906 ( .A1(n3952), .A2(n3953), .A3(n3954), .A4(n3955), .ZN(n3936)
         );
  NOR4_X2 U1907 ( .A1(u4_N6066), .A2(u4_N6065), .A3(u4_N6064), .A4(u4_N6063), 
        .ZN(n3955) );
  NOR4_X2 U1909 ( .A1(u4_N6059), .A2(u4_N6058), .A3(u4_N6057), .A4(u4_N6056), 
        .ZN(n3953) );
  AOI22_X2 U1911 ( .A1(u4_N5959), .A2(n4580), .B1(u4_N6067), .B2(n3894), .ZN(
        n3865) );
  INV_X4 U1912 ( .A(n3956), .ZN(n3894) );
  OAI211_X2 U1913 ( .C1(n3957), .C2(n2434), .A(n3958), .B(n3959), .ZN(n3956)
         );
  OAI22_X2 U1915 ( .A1(n2506), .A2(n2507), .B1(n2508), .B2(n3962), .ZN(n2485)
         );
  NAND2_X2 U1916 ( .A1(n2511), .A2(n2514), .ZN(n3962) );
  NAND2_X2 U1917 ( .A1(u4_N6463), .A2(n3545), .ZN(n2511) );
  NAND2_X2 U1918 ( .A1(n6317), .A2(n3963), .ZN(n3545) );
  NAND2_X2 U1922 ( .A1(n6095), .A2(u4_N6463), .ZN(n3476) );
  NAND2_X2 U1924 ( .A1(u4_exp_in_pl1_11_), .A2(fract_denorm[105]), .ZN(n3964)
         );
  OR2_X2 U1925 ( .A1(u4_exp_in_pl1_9_), .A2(u4_exp_in_pl1_10_), .ZN(n3961) );
  OR2_X2 U1926 ( .A1(u4_div_scht1a[10]), .A2(u4_div_scht1a[9]), .ZN(n3960) );
  AOI22_X2 U1928 ( .A1(n3489), .A2(n6448), .B1(n4356), .B2(n3533), .ZN(n2515)
         );
  NOR2_X4 U1929 ( .A1(n6447), .A2(u4_N6463), .ZN(n3533) );
  INV_X4 U1932 ( .A(u4_N6463), .ZN(n3489) );
  AOI22_X2 U1934 ( .A1(opas_r2), .A2(u4_N5837), .B1(n3843), .B2(u4_N5836), 
        .ZN(n3548) );
  NAND4_X2 U1935 ( .A1(rmode_r3[1]), .A2(rmode_r3[0]), .A3(opas_r2), .A4(n6337), .ZN(n3843) );
  AOI221_X2 U1937 ( .B1(n4575), .B2(quo[2]), .C1(n4569), .C2(prod[0]), .A(
        n3967), .ZN(n3877) );
  AND2_X2 U1938 ( .A1(fract_i2f[0]), .A2(n4662), .ZN(n3967) );
  AND3_X2 U1940 ( .A1(n3873), .A2(n2763), .A3(n2700), .ZN(n2630) );
  AND3_X2 U1941 ( .A1(n3171), .A2(n2751), .A3(n2659), .ZN(n2700) );
  NAND4_X2 U1943 ( .A1(n3968), .A2(n3969), .A3(n3970), .A4(n3971), .ZN(n2684)
         );
  NOR4_X2 U1944 ( .A1(n6444), .A2(fract_denorm[51]), .A3(fract_denorm[50]), 
        .A4(n6445), .ZN(n3971) );
  AOI221_X2 U1945 ( .B1(n4571), .B2(quo[44]), .C1(n4569), .C2(prod[42]), .A(
        n3972), .ZN(n2770) );
  AND2_X2 U1946 ( .A1(fract_i2f[42]), .A2(n4662), .ZN(n3972) );
  OAI211_X2 U1947 ( .C1(n3973), .C2(n4434), .A(n3974), .B(n3975), .ZN(
        fract_denorm[50]) );
  AOI22_X2 U1948 ( .A1(fract_out_q[1]), .A2(n4595), .B1(fract_i2f[50]), .B2(
        n4661), .ZN(n3975) );
  AOI22_X2 U1949 ( .A1(quo[0]), .A2(n4563), .B1(quo[52]), .B2(n4572), .ZN(
        n3974) );
  OAI211_X2 U1950 ( .C1(n3973), .C2(n4432), .A(n3977), .B(n3978), .ZN(
        fract_denorm[51]) );
  AOI22_X2 U1951 ( .A1(fract_out_q[2]), .A2(n4595), .B1(fract_i2f[51]), .B2(
        n4661), .ZN(n3978) );
  AOI221_X2 U1953 ( .B1(n4571), .B2(quo[11]), .C1(n4569), .C2(prod[9]), .A(
        n3979), .ZN(n2718) );
  AND2_X2 U1954 ( .A1(fract_i2f[9]), .A2(n4662), .ZN(n3979) );
  NOR4_X2 U1955 ( .A1(n6440), .A2(n6441), .A3(n6442), .A4(n6443), .ZN(n3970)
         );
  AOI221_X2 U1956 ( .B1(n4571), .B2(quo[12]), .C1(n4569), .C2(prod[10]), .A(
        n3980), .ZN(n3876) );
  AND2_X2 U1957 ( .A1(fract_i2f[10]), .A2(n4662), .ZN(n3980) );
  AOI221_X2 U1958 ( .B1(n4571), .B2(quo[20]), .C1(n4569), .C2(prod[18]), .A(
        n3981), .ZN(n2636) );
  AND2_X2 U1959 ( .A1(fract_i2f[18]), .A2(n4662), .ZN(n3981) );
  AOI221_X2 U1960 ( .B1(n4571), .B2(quo[28]), .C1(n4569), .C2(prod[26]), .A(
        n3982), .ZN(n2605) );
  AND2_X2 U1961 ( .A1(fract_i2f[26]), .A2(n4662), .ZN(n3982) );
  AOI221_X2 U1962 ( .B1(n4571), .B2(quo[36]), .C1(n4569), .C2(prod[34]), .A(
        n3983), .ZN(n2633) );
  AND2_X2 U1963 ( .A1(fract_i2f[34]), .A2(n4662), .ZN(n3983) );
  NOR4_X2 U1964 ( .A1(n2561), .A2(n2635), .A3(n2604), .A4(n2634), .ZN(n3969)
         );
  OR3_X2 U1965 ( .A1(n6433), .A2(n6434), .A3(n2697), .ZN(n2634) );
  AOI221_X2 U1968 ( .B1(n4571), .B2(quo[41]), .C1(n4569), .C2(prod[39]), .A(
        n3985), .ZN(n3984) );
  AND2_X2 U1969 ( .A1(fract_i2f[39]), .A2(n4662), .ZN(n3985) );
  AOI221_X2 U1970 ( .B1(n4571), .B2(quo[43]), .C1(n4568), .C2(prod[41]), .A(
        n3986), .ZN(n2768) );
  AND2_X2 U1971 ( .A1(fract_i2f[41]), .A2(n4662), .ZN(n3986) );
  AOI221_X2 U1972 ( .B1(n4571), .B2(quo[42]), .C1(n4568), .C2(prod[40]), .A(
        n3987), .ZN(n2680) );
  AND2_X2 U1973 ( .A1(fract_i2f[40]), .A2(n4662), .ZN(n3987) );
  AOI221_X2 U1974 ( .B1(n4571), .B2(quo[40]), .C1(n4568), .C2(prod[38]), .A(
        n3988), .ZN(n2752) );
  AND2_X2 U1975 ( .A1(fract_i2f[38]), .A2(n4662), .ZN(n3988) );
  AOI221_X2 U1976 ( .B1(n4575), .B2(quo[39]), .C1(n4568), .C2(prod[37]), .A(
        n3989), .ZN(n3174) );
  AND2_X2 U1977 ( .A1(fract_i2f[37]), .A2(n4662), .ZN(n3989) );
  AOI221_X2 U1978 ( .B1(n4575), .B2(quo[38]), .C1(n4568), .C2(prod[36]), .A(
        n3990), .ZN(n2696) );
  AND2_X2 U1979 ( .A1(fract_i2f[36]), .A2(n4662), .ZN(n3990) );
  AOI221_X2 U1980 ( .B1(n4575), .B2(quo[37]), .C1(n4568), .C2(prod[35]), .A(
        n3991), .ZN(n2758) );
  AND2_X2 U1981 ( .A1(fract_i2f[35]), .A2(n4662), .ZN(n3991) );
  AND3_X2 U1983 ( .A1(n3175), .A2(n2739), .A3(n2669), .ZN(n2708) );
  AOI221_X2 U1985 ( .B1(n4575), .B2(quo[33]), .C1(n4568), .C2(prod[31]), .A(
        n3993), .ZN(n3992) );
  AND2_X2 U1986 ( .A1(fract_i2f[31]), .A2(n4662), .ZN(n3993) );
  AOI221_X2 U1987 ( .B1(n4575), .B2(quo[35]), .C1(n4568), .C2(prod[33]), .A(
        n3994), .ZN(n2722) );
  AND2_X2 U1988 ( .A1(fract_i2f[33]), .A2(n4662), .ZN(n3994) );
  AOI221_X2 U1989 ( .B1(n4575), .B2(quo[34]), .C1(n4568), .C2(prod[32]), .A(
        n3995), .ZN(n2681) );
  AND2_X2 U1990 ( .A1(fract_i2f[32]), .A2(n4662), .ZN(n3995) );
  AOI221_X2 U1991 ( .B1(n4575), .B2(quo[32]), .C1(n4568), .C2(prod[30]), .A(
        n3996), .ZN(n2739) );
  AND2_X2 U1992 ( .A1(fract_i2f[30]), .A2(n4662), .ZN(n3996) );
  AOI221_X2 U1993 ( .B1(n4575), .B2(quo[31]), .C1(n4568), .C2(prod[29]), .A(
        n3997), .ZN(n3175) );
  AND2_X2 U1994 ( .A1(fract_i2f[29]), .A2(n4662), .ZN(n3997) );
  AOI221_X2 U1995 ( .B1(n4575), .B2(quo[30]), .C1(n4568), .C2(prod[28]), .A(
        n3998), .ZN(n2730) );
  AND2_X2 U1996 ( .A1(fract_i2f[28]), .A2(n4662), .ZN(n3998) );
  AOI221_X2 U1997 ( .B1(n4575), .B2(quo[29]), .C1(n4568), .C2(prod[27]), .A(
        n3999), .ZN(n3176) );
  AND2_X2 U1998 ( .A1(fract_i2f[27]), .A2(n4662), .ZN(n3999) );
  AND3_X2 U2000 ( .A1(n3177), .A2(n2753), .A3(n2660), .ZN(n2695) );
  AOI221_X2 U2002 ( .B1(n4575), .B2(quo[25]), .C1(n4568), .C2(prod[23]), .A(
        n4001), .ZN(n4000) );
  AND2_X2 U2003 ( .A1(fract_i2f[23]), .A2(n4662), .ZN(n4001) );
  AOI221_X2 U2004 ( .B1(n4572), .B2(quo[27]), .C1(n4568), .C2(prod[25]), .A(
        n4002), .ZN(n2685) );
  AND2_X2 U2005 ( .A1(fract_i2f[25]), .A2(n4662), .ZN(n4002) );
  AOI221_X2 U2006 ( .B1(n4572), .B2(quo[26]), .C1(n4568), .C2(prod[24]), .A(
        n4003), .ZN(n2769) );
  AND2_X2 U2007 ( .A1(fract_i2f[24]), .A2(n4662), .ZN(n4003) );
  AOI221_X2 U2008 ( .B1(n4572), .B2(quo[24]), .C1(n4568), .C2(prod[22]), .A(
        n4004), .ZN(n2753) );
  AND2_X2 U2009 ( .A1(fract_i2f[22]), .A2(n4662), .ZN(n4004) );
  AOI221_X2 U2010 ( .B1(n4572), .B2(quo[23]), .C1(n4568), .C2(prod[21]), .A(
        n4005), .ZN(n3177) );
  AND2_X2 U2011 ( .A1(fract_i2f[21]), .A2(n4662), .ZN(n4005) );
  AOI221_X2 U2012 ( .B1(n4572), .B2(quo[22]), .C1(n4568), .C2(prod[20]), .A(
        n4006), .ZN(n2762) );
  AND2_X2 U2013 ( .A1(fract_i2f[20]), .A2(n4662), .ZN(n4006) );
  AOI221_X2 U2014 ( .B1(n4572), .B2(quo[21]), .C1(n4568), .C2(prod[19]), .A(
        n4007), .ZN(n3178) );
  AND2_X2 U2015 ( .A1(fract_i2f[19]), .A2(n4662), .ZN(n4007) );
  AND3_X2 U2017 ( .A1(n3179), .A2(n2740), .A3(n2670), .ZN(n2709) );
  AOI221_X2 U2019 ( .B1(n4572), .B2(quo[17]), .C1(n4568), .C2(prod[15]), .A(
        n4009), .ZN(n4008) );
  AND2_X2 U2020 ( .A1(fract_i2f[15]), .A2(n4662), .ZN(n4009) );
  AOI221_X2 U2021 ( .B1(n4572), .B2(quo[19]), .C1(n4568), .C2(prod[17]), .A(
        n4010), .ZN(n2593) );
  AND2_X2 U2022 ( .A1(fract_i2f[17]), .A2(n4662), .ZN(n4010) );
  AOI221_X2 U2023 ( .B1(n4572), .B2(quo[18]), .C1(n4568), .C2(prod[16]), .A(
        n4011), .ZN(n2745) );
  AND2_X2 U2024 ( .A1(fract_i2f[16]), .A2(n4662), .ZN(n4011) );
  AOI221_X2 U2025 ( .B1(n4572), .B2(quo[16]), .C1(n4568), .C2(prod[14]), .A(
        n4012), .ZN(n2740) );
  AND2_X2 U2026 ( .A1(fract_i2f[14]), .A2(n4662), .ZN(n4012) );
  AOI221_X2 U2027 ( .B1(n4572), .B2(quo[15]), .C1(n4568), .C2(prod[13]), .A(
        n4013), .ZN(n3179) );
  AND2_X2 U2028 ( .A1(fract_i2f[13]), .A2(n4662), .ZN(n4013) );
  AOI221_X2 U2029 ( .B1(n4574), .B2(quo[14]), .C1(n4568), .C2(prod[12]), .A(
        n4014), .ZN(n2731) );
  AND2_X2 U2030 ( .A1(fract_i2f[12]), .A2(n4662), .ZN(n4014) );
  AOI221_X2 U2031 ( .B1(n4572), .B2(quo[13]), .C1(n4568), .C2(prod[11]), .A(
        n4015), .ZN(n3180) );
  AND2_X2 U2032 ( .A1(fract_i2f[11]), .A2(fpu_op_r3[2]), .ZN(n4015) );
  NAND4_X2 U2034 ( .A1(n2698), .A2(n2644), .A3(n4016), .A4(n4017), .ZN(n3912)
         );
  NOR4_X2 U2035 ( .A1(n4018), .A2(fract_denorm[66]), .A3(fract_denorm[82]), 
        .A4(fract_denorm[74]), .ZN(n4017) );
  OAI211_X2 U2036 ( .C1(n3973), .C2(n4298), .A(n4019), .B(n4020), .ZN(
        fract_denorm[74]) );
  AOI22_X2 U2037 ( .A1(fract_out_q[25]), .A2(n4595), .B1(fract_i2f[74]), .B2(
        n4661), .ZN(n4020) );
  AOI22_X2 U2038 ( .A1(quo[24]), .A2(n4563), .B1(quo[76]), .B2(n4575), .ZN(
        n4019) );
  OAI211_X2 U2039 ( .C1(n3973), .C2(n4416), .A(n4021), .B(n4022), .ZN(
        fract_denorm[82]) );
  AOI22_X2 U2040 ( .A1(fract_out_q[33]), .A2(n4595), .B1(fract_i2f[82]), .B2(
        n4661), .ZN(n4022) );
  AOI22_X2 U2041 ( .A1(quo[32]), .A2(n4563), .B1(quo[84]), .B2(n4575), .ZN(
        n4021) );
  OAI211_X2 U2042 ( .C1(n3973), .C2(n4423), .A(n4023), .B(n4024), .ZN(
        fract_denorm[66]) );
  AOI22_X2 U2043 ( .A1(fract_out_q[17]), .A2(n4595), .B1(fract_i2f[66]), .B2(
        n4661), .ZN(n4024) );
  AOI22_X2 U2044 ( .A1(quo[16]), .A2(n4563), .B1(quo[68]), .B2(n4574), .ZN(
        n4023) );
  NAND2_X2 U2045 ( .A1(n6400), .A2(n6401), .ZN(n4018) );
  OAI211_X2 U2046 ( .C1(n3973), .C2(n4430), .A(n4025), .B(n4026), .ZN(
        fract_denorm[58]) );
  AOI22_X2 U2047 ( .A1(fract_out_q[9]), .A2(n4595), .B1(fract_i2f[58]), .B2(
        n4661), .ZN(n4026) );
  AOI22_X2 U2048 ( .A1(quo[8]), .A2(n4563), .B1(quo[60]), .B2(n4575), .ZN(
        n4025) );
  OAI211_X2 U2049 ( .C1(n3973), .C2(n4429), .A(n4027), .B(n4028), .ZN(
        fract_denorm[52]) );
  AOI22_X2 U2050 ( .A1(fract_out_q[3]), .A2(n4595), .B1(fract_i2f[52]), .B2(
        n4661), .ZN(n4028) );
  OAI211_X2 U2056 ( .C1(n3973), .C2(n4422), .A(n4029), .B(n4030), .ZN(
        fract_denorm[71]) );
  AOI22_X2 U2057 ( .A1(fract_out_q[22]), .A2(n4595), .B1(fract_i2f[71]), .B2(
        n4661), .ZN(n4030) );
  AOI22_X2 U2058 ( .A1(quo[21]), .A2(n4563), .B1(quo[73]), .B2(n4571), .ZN(
        n4029) );
  OAI211_X2 U2059 ( .C1(n3973), .C2(n4407), .A(n4031), .B(n4032), .ZN(
        fract_denorm[73]) );
  AOI22_X2 U2060 ( .A1(fract_out_q[24]), .A2(n4595), .B1(fract_i2f[73]), .B2(
        n4661), .ZN(n4032) );
  AOI22_X2 U2061 ( .A1(quo[23]), .A2(n4563), .B1(quo[75]), .B2(n4574), .ZN(
        n4031) );
  OAI211_X2 U2062 ( .C1(n3973), .C2(n4313), .A(n4033), .B(n4034), .ZN(
        fract_denorm[72]) );
  AOI22_X2 U2063 ( .A1(fract_out_q[23]), .A2(n4595), .B1(fract_i2f[72]), .B2(
        n4661), .ZN(n4034) );
  AOI22_X2 U2064 ( .A1(quo[22]), .A2(n4563), .B1(quo[74]), .B2(n4575), .ZN(
        n4033) );
  OAI211_X2 U2065 ( .C1(n3973), .C2(n4415), .A(n4035), .B(n4036), .ZN(
        fract_denorm[70]) );
  AOI22_X2 U2066 ( .A1(fract_out_q[21]), .A2(n4595), .B1(fract_i2f[70]), .B2(
        n4661), .ZN(n4036) );
  AOI22_X2 U2067 ( .A1(quo[20]), .A2(n4563), .B1(quo[72]), .B2(n4574), .ZN(
        n4035) );
  OAI211_X2 U2068 ( .C1(n4567), .C2(n4342), .A(n4037), .B(n4038), .ZN(
        fract_denorm[69]) );
  AOI22_X2 U2069 ( .A1(fract_out_q[20]), .A2(n4595), .B1(fract_i2f[69]), .B2(
        n4661), .ZN(n4038) );
  AOI22_X2 U2070 ( .A1(quo[19]), .A2(n4563), .B1(quo[71]), .B2(n4574), .ZN(
        n4037) );
  OAI211_X2 U2071 ( .C1(n4567), .C2(n4402), .A(n4039), .B(n4040), .ZN(
        fract_denorm[68]) );
  AOI22_X2 U2072 ( .A1(fract_out_q[19]), .A2(n4595), .B1(fract_i2f[68]), .B2(
        n4661), .ZN(n4040) );
  AOI22_X2 U2073 ( .A1(quo[18]), .A2(n4563), .B1(quo[70]), .B2(n4574), .ZN(
        n4039) );
  OAI211_X2 U2074 ( .C1(n4567), .C2(n4311), .A(n4041), .B(n4042), .ZN(
        fract_denorm[67]) );
  AOI22_X2 U2075 ( .A1(fract_out_q[18]), .A2(n4595), .B1(fract_i2f[67]), .B2(
        n4661), .ZN(n4042) );
  AOI22_X2 U2076 ( .A1(quo[17]), .A2(n4563), .B1(quo[69]), .B2(n4575), .ZN(
        n4041) );
  OR3_X2 U2077 ( .A1(fract_denorm[59]), .A2(fract_denorm[60]), .A3(n6388), 
        .ZN(n2592) );
  OAI211_X2 U2080 ( .C1(n4567), .C2(n4297), .A(n4043), .B(n4044), .ZN(
        fract_denorm[63]) );
  AOI22_X2 U2081 ( .A1(fract_out_q[14]), .A2(n4595), .B1(fract_i2f[63]), .B2(
        n4661), .ZN(n4044) );
  AOI22_X2 U2082 ( .A1(quo[13]), .A2(n4563), .B1(quo[65]), .B2(n4574), .ZN(
        n4043) );
  OAI211_X2 U2083 ( .C1(n4567), .C2(n4414), .A(n4045), .B(n4046), .ZN(
        fract_denorm[65]) );
  AOI22_X2 U2084 ( .A1(fract_out_q[16]), .A2(n4595), .B1(fract_i2f[65]), .B2(
        n4662), .ZN(n4046) );
  AOI22_X2 U2085 ( .A1(quo[15]), .A2(n4563), .B1(quo[67]), .B2(n4574), .ZN(
        n4045) );
  OAI211_X2 U2086 ( .C1(n4567), .C2(n4428), .A(n4047), .B(n4048), .ZN(
        fract_denorm[64]) );
  AOI22_X2 U2087 ( .A1(fract_out_q[15]), .A2(n4595), .B1(fract_i2f[64]), .B2(
        n4662), .ZN(n4048) );
  AOI22_X2 U2088 ( .A1(quo[14]), .A2(n4563), .B1(quo[66]), .B2(n4574), .ZN(
        n4047) );
  OAI211_X2 U2089 ( .C1(n4567), .C2(n4312), .A(n4049), .B(n4050), .ZN(
        fract_denorm[62]) );
  AOI22_X2 U2090 ( .A1(fract_out_q[13]), .A2(n4595), .B1(fract_i2f[62]), .B2(
        n4662), .ZN(n4050) );
  AOI22_X2 U2091 ( .A1(quo[12]), .A2(n4563), .B1(quo[64]), .B2(n4574), .ZN(
        n4049) );
  OAI211_X2 U2092 ( .C1(n4567), .C2(n4406), .A(n4051), .B(n4052), .ZN(
        fract_denorm[61]) );
  AOI22_X2 U2093 ( .A1(fract_out_q[12]), .A2(n4595), .B1(fract_i2f[61]), .B2(
        n4662), .ZN(n4052) );
  AOI22_X2 U2094 ( .A1(quo[11]), .A2(n4563), .B1(quo[63]), .B2(n4573), .ZN(
        n4051) );
  OAI211_X2 U2095 ( .C1(n4567), .C2(n4346), .A(n4053), .B(n4054), .ZN(
        fract_denorm[60]) );
  AOI22_X2 U2096 ( .A1(fract_out_q[11]), .A2(n4595), .B1(fract_i2f[60]), .B2(
        n4662), .ZN(n4054) );
  AOI22_X2 U2097 ( .A1(quo[10]), .A2(n4563), .B1(quo[62]), .B2(n4575), .ZN(
        n4053) );
  OAI211_X2 U2098 ( .C1(n4567), .C2(n4413), .A(n4055), .B(n4056), .ZN(
        fract_denorm[59]) );
  AOI22_X2 U2099 ( .A1(fract_out_q[10]), .A2(n4595), .B1(fract_i2f[59]), .B2(
        n4662), .ZN(n4056) );
  AOI22_X2 U2100 ( .A1(quo[9]), .A2(n4563), .B1(quo[61]), .B2(n4573), .ZN(
        n4055) );
  OAI211_X2 U2104 ( .C1(n4567), .C2(n4436), .A(n4057), .B(n4058), .ZN(
        fract_denorm[79]) );
  AOI22_X2 U2105 ( .A1(fract_out_q[30]), .A2(n4595), .B1(fract_i2f[79]), .B2(
        n4662), .ZN(n4058) );
  AOI22_X2 U2106 ( .A1(quo[29]), .A2(n4563), .B1(quo[81]), .B2(n4571), .ZN(
        n4057) );
  OAI211_X2 U2107 ( .C1(n4566), .C2(n4427), .A(n4059), .B(n4060), .ZN(
        fract_denorm[81]) );
  AOI22_X2 U2108 ( .A1(fract_out_q[32]), .A2(n4595), .B1(fract_i2f[81]), .B2(
        n4662), .ZN(n4060) );
  AOI22_X2 U2109 ( .A1(quo[31]), .A2(n4563), .B1(quo[83]), .B2(n4573), .ZN(
        n4059) );
  OAI211_X2 U2110 ( .C1(n4566), .C2(n4437), .A(n4061), .B(n4062), .ZN(
        fract_denorm[80]) );
  AOI22_X2 U2111 ( .A1(fract_out_q[31]), .A2(n4595), .B1(fract_i2f[80]), .B2(
        n4662), .ZN(n4062) );
  AOI22_X2 U2112 ( .A1(quo[30]), .A2(n4563), .B1(quo[82]), .B2(n4574), .ZN(
        n4061) );
  OAI211_X2 U2113 ( .C1(n4566), .C2(n4421), .A(n4063), .B(n4064), .ZN(
        fract_denorm[78]) );
  AOI22_X2 U2114 ( .A1(fract_out_q[29]), .A2(n4595), .B1(fract_i2f[78]), .B2(
        n4662), .ZN(n4064) );
  AOI22_X2 U2115 ( .A1(quo[28]), .A2(n4563), .B1(quo[80]), .B2(n4573), .ZN(
        n4063) );
  OAI211_X2 U2116 ( .C1(n3973), .C2(n4412), .A(n4065), .B(n4066), .ZN(
        fract_denorm[77]) );
  AOI22_X2 U2117 ( .A1(fract_out_q[28]), .A2(n4595), .B1(fract_i2f[77]), .B2(
        n4662), .ZN(n4066) );
  AOI22_X2 U2118 ( .A1(quo[27]), .A2(n4563), .B1(quo[79]), .B2(n4575), .ZN(
        n4065) );
  OAI211_X2 U2119 ( .C1(n3973), .C2(n4426), .A(n4067), .B(n4068), .ZN(
        fract_denorm[76]) );
  AOI22_X2 U2120 ( .A1(fract_out_q[27]), .A2(n4595), .B1(fract_i2f[76]), .B2(
        n4662), .ZN(n4068) );
  AOI22_X2 U2121 ( .A1(quo[26]), .A2(n4563), .B1(quo[78]), .B2(n4573), .ZN(
        n4067) );
  OAI211_X2 U2122 ( .C1(n3973), .C2(n4343), .A(n4069), .B(n4070), .ZN(
        fract_denorm[75]) );
  AOI22_X2 U2123 ( .A1(fract_out_q[26]), .A2(n4595), .B1(fract_i2f[75]), .B2(
        n4662), .ZN(n4070) );
  AOI22_X2 U2124 ( .A1(quo[25]), .A2(n4563), .B1(quo[77]), .B2(n4575), .ZN(
        n4069) );
  OAI211_X2 U2128 ( .C1(n3973), .C2(n4294), .A(n4071), .B(n4072), .ZN(
        fract_denorm[87]) );
  AOI22_X2 U2129 ( .A1(fract_out_q[38]), .A2(n4595), .B1(fract_i2f[87]), .B2(
        n4662), .ZN(n4072) );
  AOI22_X2 U2130 ( .A1(quo[37]), .A2(n4563), .B1(quo[89]), .B2(n4571), .ZN(
        n4071) );
  OAI211_X2 U2131 ( .C1(n3973), .C2(n4411), .A(n4073), .B(n4074), .ZN(
        fract_denorm[89]) );
  AOI22_X2 U2132 ( .A1(fract_out_q[40]), .A2(n4595), .B1(fract_i2f[89]), .B2(
        n4662), .ZN(n4074) );
  AOI22_X2 U2133 ( .A1(quo[39]), .A2(n4563), .B1(quo[91]), .B2(n4574), .ZN(
        n4073) );
  OAI211_X2 U2134 ( .C1(n3973), .C2(n4425), .A(n4075), .B(n4076), .ZN(
        fract_denorm[88]) );
  AOI22_X2 U2135 ( .A1(fract_out_q[39]), .A2(n4595), .B1(fract_i2f[88]), .B2(
        n4662), .ZN(n4076) );
  AOI22_X2 U2136 ( .A1(quo[38]), .A2(n4563), .B1(quo[90]), .B2(n4572), .ZN(
        n4075) );
  OAI211_X2 U2137 ( .C1(n3973), .C2(n4307), .A(n4077), .B(n4078), .ZN(
        fract_denorm[86]) );
  AOI22_X2 U2138 ( .A1(fract_out_q[37]), .A2(n4595), .B1(fract_i2f[86]), .B2(
        n4662), .ZN(n4078) );
  AOI22_X2 U2139 ( .A1(quo[36]), .A2(n4563), .B1(quo[88]), .B2(n4574), .ZN(
        n4077) );
  OAI211_X2 U2140 ( .C1(n3973), .C2(n4404), .A(n4079), .B(n4080), .ZN(
        fract_denorm[85]) );
  AOI22_X2 U2141 ( .A1(fract_out_q[36]), .A2(n4595), .B1(fract_i2f[85]), .B2(
        n4662), .ZN(n4080) );
  AOI22_X2 U2142 ( .A1(quo[35]), .A2(n4563), .B1(quo[87]), .B2(n4571), .ZN(
        n4079) );
  OAI211_X2 U2143 ( .C1(n4567), .C2(n4344), .A(n4081), .B(n4082), .ZN(
        fract_denorm[84]) );
  AOI22_X2 U2144 ( .A1(fract_out_q[35]), .A2(n4595), .B1(fract_i2f[84]), .B2(
        n4662), .ZN(n4082) );
  AOI22_X2 U2145 ( .A1(quo[34]), .A2(n4564), .B1(quo[86]), .B2(n4573), .ZN(
        n4081) );
  OAI211_X2 U2146 ( .C1(n4567), .C2(n4420), .A(n4083), .B(n4084), .ZN(
        fract_denorm[83]) );
  AOI22_X2 U2147 ( .A1(fract_out_q[34]), .A2(n4595), .B1(fract_i2f[83]), .B2(
        n4662), .ZN(n4084) );
  AOI22_X2 U2148 ( .A1(quo[33]), .A2(n4564), .B1(quo[85]), .B2(n4571), .ZN(
        n4083) );
  OAI211_X2 U2151 ( .C1(n4567), .C2(n4310), .A(n4085), .B(n4086), .ZN(
        fract_denorm[55]) );
  AOI22_X2 U2152 ( .A1(fract_out_q[6]), .A2(n4595), .B1(fract_i2f[55]), .B2(
        n4662), .ZN(n4086) );
  AOI22_X2 U2153 ( .A1(quo[5]), .A2(n4564), .B1(quo[57]), .B2(n4575), .ZN(
        n4085) );
  OAI211_X2 U2154 ( .C1(n4567), .C2(n4341), .A(n4087), .B(n4088), .ZN(
        fract_denorm[57]) );
  AOI22_X2 U2155 ( .A1(fract_out_q[8]), .A2(n4595), .B1(fract_i2f[57]), .B2(
        n4662), .ZN(n4088) );
  AOI22_X2 U2156 ( .A1(quo[7]), .A2(n4564), .B1(quo[59]), .B2(n4575), .ZN(
        n4087) );
  OAI211_X2 U2157 ( .C1(n4567), .C2(n4401), .A(n4089), .B(n4090), .ZN(
        fract_denorm[56]) );
  AOI22_X2 U2158 ( .A1(fract_out_q[7]), .A2(n4595), .B1(fract_i2f[56]), .B2(
        n4662), .ZN(n4090) );
  AOI22_X2 U2159 ( .A1(quo[6]), .A2(n4564), .B1(quo[58]), .B2(n4575), .ZN(
        n4089) );
  OAI211_X2 U2160 ( .C1(n4567), .C2(n4419), .A(n4091), .B(n4092), .ZN(
        fract_denorm[54]) );
  AOI22_X2 U2161 ( .A1(fract_out_q[5]), .A2(n4595), .B1(fract_i2f[54]), .B2(
        n4662), .ZN(n4092) );
  AOI22_X2 U2162 ( .A1(quo[4]), .A2(n4564), .B1(quo[56]), .B2(n4575), .ZN(
        n4091) );
  OAI211_X2 U2163 ( .C1(n4567), .C2(n4410), .A(n4093), .B(n4094), .ZN(
        fract_denorm[53]) );
  AOI22_X2 U2164 ( .A1(fract_out_q[4]), .A2(n4595), .B1(fract_i2f[53]), .B2(
        fpu_op_r3[2]), .ZN(n4094) );
  AOI22_X2 U2165 ( .A1(quo[3]), .A2(n4564), .B1(quo[55]), .B2(n4571), .ZN(
        n4093) );
  AND3_X2 U2167 ( .A1(n3172), .A2(n2737), .A3(n2668), .ZN(n2706) );
  AOI221_X2 U2169 ( .B1(n4571), .B2(quo[49]), .C1(n4568), .C2(prod[47]), .A(
        n4096), .ZN(n4095) );
  AND2_X2 U2170 ( .A1(fract_i2f[47]), .A2(fpu_op_r3[2]), .ZN(n4096) );
  AOI221_X2 U2171 ( .B1(n4573), .B2(quo[51]), .C1(n4568), .C2(prod[49]), .A(
        n6368), .ZN(n2711) );
  AOI22_X2 U2172 ( .A1(fract_out_q[0]), .A2(n4595), .B1(fract_i2f[49]), .B2(
        fpu_op_r3[2]), .ZN(n4097) );
  AOI221_X2 U2173 ( .B1(n4573), .B2(quo[50]), .C1(n4568), .C2(prod[48]), .A(
        n4098), .ZN(n2744) );
  AND2_X2 U2174 ( .A1(fract_i2f[48]), .A2(fpu_op_r3[2]), .ZN(n4098) );
  AOI221_X2 U2175 ( .B1(n4573), .B2(quo[48]), .C1(n4568), .C2(prod[46]), .A(
        n4099), .ZN(n2737) );
  AND2_X2 U2176 ( .A1(fract_i2f[46]), .A2(fpu_op_r3[2]), .ZN(n4099) );
  AOI221_X2 U2177 ( .B1(n4571), .B2(quo[47]), .C1(n4568), .C2(prod[45]), .A(
        n4100), .ZN(n3172) );
  AND2_X2 U2178 ( .A1(fract_i2f[45]), .A2(fpu_op_r3[2]), .ZN(n4100) );
  AOI221_X2 U2179 ( .B1(n4573), .B2(quo[46]), .C1(n4568), .C2(prod[44]), .A(
        n4101), .ZN(n2729) );
  AND2_X2 U2180 ( .A1(fract_i2f[44]), .A2(fpu_op_r3[2]), .ZN(n4101) );
  AOI221_X2 U2181 ( .B1(n4573), .B2(quo[45]), .C1(n4568), .C2(prod[43]), .A(
        n4102), .ZN(n3173) );
  AND2_X2 U2182 ( .A1(fract_i2f[43]), .A2(fpu_op_r3[2]), .ZN(n4102) );
  NAND2_X2 U2184 ( .A1(n2638), .A2(n6365), .ZN(n2598) );
  OAI211_X2 U2185 ( .C1(n4566), .C2(n4435), .A(n4103), .B(n4104), .ZN(
        fract_denorm[98]) );
  AOI22_X2 U2186 ( .A1(fract_out_q[49]), .A2(n3315), .B1(fract_i2f[98]), .B2(
        n4661), .ZN(n4104) );
  AOI22_X2 U2187 ( .A1(quo[48]), .A2(n4564), .B1(quo[100]), .B2(n4571), .ZN(
        n4103) );
  AND3_X2 U2188 ( .A1(n6360), .A2(n4654), .A3(n2761), .ZN(n2638) );
  OR3_X2 U2190 ( .A1(fract_denorm[101]), .A2(fract_denorm[102]), .A3(
        fract_denorm[100]), .ZN(n2662) );
  OAI211_X2 U2191 ( .C1(n4566), .C2(n4409), .A(n4105), .B(n4106), .ZN(
        fract_denorm[100]) );
  AOI22_X2 U2192 ( .A1(fract_out_q[51]), .A2(n3315), .B1(fract_i2f[100]), .B2(
        n4661), .ZN(n4106) );
  AOI22_X2 U2193 ( .A1(quo[50]), .A2(n4309), .B1(quo[102]), .B2(n4570), .ZN(
        n4105) );
  OAI211_X2 U2194 ( .C1(n4566), .C2(n4306), .A(n4107), .B(n4108), .ZN(
        fract_denorm[102]) );
  AOI22_X2 U2195 ( .A1(fract_out_q[53]), .A2(n3315), .B1(fract_i2f[102]), .B2(
        n4661), .ZN(n4108) );
  AOI22_X2 U2196 ( .A1(quo[52]), .A2(n4309), .B1(quo[104]), .B2(n4570), .ZN(
        n4107) );
  OAI211_X2 U2197 ( .C1(n4566), .C2(n4418), .A(n4109), .B(n4110), .ZN(
        fract_denorm[101]) );
  AOI22_X2 U2198 ( .A1(fract_out_q[52]), .A2(n3315), .B1(fract_i2f[101]), .B2(
        n4662), .ZN(n4110) );
  AOI22_X2 U2199 ( .A1(quo[51]), .A2(n4309), .B1(quo[103]), .B2(n4570), .ZN(
        n4109) );
  OAI211_X2 U2200 ( .C1(n4566), .C2(n4338), .A(n4111), .B(n4112), .ZN(
        fract_denorm[104]) );
  AOI22_X2 U2201 ( .A1(fract_out_q[55]), .A2(n3315), .B1(fract_i2f[104]), .B2(
        n4661), .ZN(n4112) );
  OAI211_X2 U2203 ( .C1(n4566), .C2(n4403), .A(n4113), .B(n4114), .ZN(
        fract_denorm[103]) );
  AOI22_X2 U2204 ( .A1(fract_out_q[54]), .A2(n3315), .B1(fract_i2f[103]), .B2(
        n4661), .ZN(n4114) );
  OAI211_X2 U2206 ( .C1(n4566), .C2(n4433), .A(n4115), .B(n4116), .ZN(
        fract_denorm[99]) );
  AOI22_X2 U2207 ( .A1(fract_out_q[50]), .A2(n4595), .B1(fract_i2f[99]), .B2(
        n4662), .ZN(n4116) );
  AOI22_X2 U2208 ( .A1(quo[49]), .A2(n4564), .B1(quo[101]), .B2(n4571), .ZN(
        n4115) );
  OAI211_X2 U2209 ( .C1(n4566), .C2(n4345), .A(n4117), .B(n4118), .ZN(
        fract_denorm[90]) );
  AOI22_X2 U2210 ( .A1(fract_out_q[41]), .A2(n3315), .B1(fract_i2f[90]), .B2(
        n4661), .ZN(n4118) );
  AOI22_X2 U2211 ( .A1(quo[40]), .A2(n4564), .B1(quo[92]), .B2(n4571), .ZN(
        n4117) );
  OAI211_X2 U2215 ( .C1(n4566), .C2(n4408), .A(n4119), .B(n4120), .ZN(
        fract_denorm[95]) );
  AOI22_X2 U2216 ( .A1(fract_out_q[46]), .A2(n3315), .B1(fract_i2f[95]), .B2(
        n4661), .ZN(n4120) );
  AOI22_X2 U2217 ( .A1(quo[45]), .A2(n4564), .B1(quo[97]), .B2(n4572), .ZN(
        n4119) );
  OAI211_X2 U2218 ( .C1(n4566), .C2(n4431), .A(n4121), .B(n4122), .ZN(
        fract_denorm[97]) );
  AOI22_X2 U2219 ( .A1(fract_out_q[48]), .A2(n3315), .B1(fract_i2f[97]), .B2(
        n4661), .ZN(n4122) );
  AOI22_X2 U2220 ( .A1(quo[47]), .A2(n4564), .B1(quo[99]), .B2(n4573), .ZN(
        n4121) );
  OAI211_X2 U2221 ( .C1(n4566), .C2(n4417), .A(n4123), .B(n4124), .ZN(
        fract_denorm[96]) );
  AOI22_X2 U2222 ( .A1(fract_out_q[47]), .A2(n4595), .B1(fract_i2f[96]), .B2(
        n4661), .ZN(n4124) );
  AOI22_X2 U2223 ( .A1(quo[46]), .A2(n4564), .B1(quo[98]), .B2(n4571), .ZN(
        n4123) );
  OAI211_X2 U2224 ( .C1(n4566), .C2(n4424), .A(n4125), .B(n4126), .ZN(
        fract_denorm[94]) );
  AOI22_X2 U2225 ( .A1(fract_out_q[45]), .A2(n3315), .B1(fract_i2f[94]), .B2(
        n4661), .ZN(n4126) );
  AOI22_X2 U2226 ( .A1(quo[44]), .A2(n4564), .B1(quo[96]), .B2(n4572), .ZN(
        n4125) );
  OAI211_X2 U2227 ( .C1(n4566), .C2(n4295), .A(n4127), .B(n4128), .ZN(
        fract_denorm[93]) );
  AOI22_X2 U2228 ( .A1(fract_out_q[44]), .A2(n3315), .B1(fract_i2f[93]), .B2(
        n4661), .ZN(n4128) );
  AOI22_X2 U2229 ( .A1(quo[43]), .A2(n4564), .B1(quo[95]), .B2(n4572), .ZN(
        n4127) );
  OAI211_X2 U2230 ( .C1(n4566), .C2(n4308), .A(n4129), .B(n4130), .ZN(
        fract_denorm[92]) );
  AOI22_X2 U2231 ( .A1(fract_out_q[43]), .A2(n3315), .B1(fract_i2f[92]), .B2(
        n4662), .ZN(n4130) );
  AOI22_X2 U2232 ( .A1(quo[42]), .A2(n4564), .B1(quo[94]), .B2(n4575), .ZN(
        n4129) );
  OAI211_X2 U2233 ( .C1(n4566), .C2(n4405), .A(n4131), .B(n4132), .ZN(
        fract_denorm[91]) );
  AOI22_X2 U2234 ( .A1(fract_out_q[42]), .A2(n4595), .B1(fract_i2f[91]), .B2(
        n4661), .ZN(n4132) );
  AOI22_X2 U2236 ( .A1(quo[41]), .A2(n4564), .B1(quo[93]), .B2(n4571), .ZN(
        n4131) );
  AOI221_X2 U2238 ( .B1(n4571), .B2(quo[10]), .C1(n4568), .C2(prod[8]), .A(
        n4133), .ZN(n2683) );
  AND2_X2 U2239 ( .A1(fract_i2f[8]), .A2(fpu_op_r3[2]), .ZN(n4133) );
  AOI221_X2 U2240 ( .B1(n4573), .B2(quo[9]), .C1(n4568), .C2(prod[7]), .A(
        n4134), .ZN(n2767) );
  AND2_X2 U2241 ( .A1(fract_i2f[7]), .A2(fpu_op_r3[2]), .ZN(n4134) );
  AOI221_X2 U2242 ( .B1(n4573), .B2(quo[8]), .C1(n4568), .C2(prod[6]), .A(
        n4135), .ZN(n2751) );
  AND2_X2 U2243 ( .A1(fract_i2f[6]), .A2(fpu_op_r3[2]), .ZN(n4135) );
  AOI221_X2 U2244 ( .B1(n4573), .B2(quo[7]), .C1(n4568), .C2(prod[5]), .A(
        n4136), .ZN(n3171) );
  AND2_X2 U2245 ( .A1(fract_i2f[5]), .A2(fpu_op_r3[2]), .ZN(n4136) );
  AOI221_X2 U2246 ( .B1(n4574), .B2(quo[6]), .C1(n4568), .C2(prod[4]), .A(
        n4137), .ZN(n2763) );
  AND2_X2 U2247 ( .A1(fract_i2f[4]), .A2(n4662), .ZN(n4137) );
  AOI221_X2 U2248 ( .B1(n4573), .B2(quo[5]), .C1(n4568), .C2(prod[3]), .A(
        n4138), .ZN(n3873) );
  AND2_X2 U2249 ( .A1(fract_i2f[3]), .A2(n4662), .ZN(n4138) );
  AOI221_X2 U2250 ( .B1(n4572), .B2(quo[4]), .C1(n4569), .C2(prod[2]), .A(
        n4139), .ZN(n2724) );
  AND2_X2 U2251 ( .A1(fract_i2f[2]), .A2(n4662), .ZN(n4139) );
  AOI221_X2 U2252 ( .B1(n4571), .B2(quo[3]), .C1(n4568), .C2(prod[1]), .A(
        n4140), .ZN(n3879) );
  AND2_X2 U2253 ( .A1(fract_i2f[1]), .A2(n4662), .ZN(n4140) );
  OAI221_X2 U2256 ( .B1(n6340), .B2(n6460), .C1(n2441), .C2(n4540), .A(n4141), 
        .ZN(n3958) );
  AND2_X2 U2258 ( .A1(n2479), .A2(n3913), .ZN(n2478) );
  NAND2_X2 U2259 ( .A1(exp_ovf_r[1]), .A2(n3488), .ZN(n3913) );
  NAND4_X2 U2265 ( .A1(n4299), .A2(n4347), .A3(n4142), .A4(n4143), .ZN(n2514)
         );
  NOR4_X2 U2266 ( .A1(n4144), .A2(exp_r[1]), .A3(n4655), .A4(n4315), .ZN(n4143) );
  NAND2_X2 U2267 ( .A1(n3965), .A2(n4349), .ZN(n4144) );
  NAND2_X2 U2270 ( .A1(n4145), .A2(n4146), .ZN(n3495) );
  NOR4_X2 U2271 ( .A1(n4147), .A2(n4148), .A3(n4149), .A4(n4150), .ZN(n4146)
         );
  NAND4_X2 U2272 ( .A1(n4151), .A2(n4152), .A3(n4153), .A4(n4154), .ZN(n4150)
         );
  NOR4_X2 U2273 ( .A1(remainder[62]), .A2(remainder[61]), .A3(remainder[60]), 
        .A4(remainder[5]), .ZN(n4154) );
  NAND4_X2 U2277 ( .A1(n4155), .A2(n4156), .A3(n4157), .A4(n4158), .ZN(n4149)
         );
  NOR4_X2 U2278 ( .A1(remainder[75]), .A2(remainder[74]), .A3(remainder[73]), 
        .A4(remainder[72]), .ZN(n4158) );
  NOR4_X2 U2280 ( .A1(remainder[69]), .A2(remainder[68]), .A3(remainder[67]), 
        .A4(remainder[66]), .ZN(n4156) );
  NAND4_X2 U2282 ( .A1(n4159), .A2(n4160), .A3(n4161), .A4(n4162), .ZN(n4148)
         );
  NOR4_X2 U2283 ( .A1(remainder[87]), .A2(remainder[86]), .A3(remainder[85]), 
        .A4(remainder[84]), .ZN(n4162) );
  NAND4_X2 U2287 ( .A1(n4163), .A2(n4164), .A3(n4165), .A4(n4166), .ZN(n4147)
         );
  NOR4_X2 U2288 ( .A1(remainder[9]), .A2(remainder[99]), .A3(remainder[98]), 
        .A4(remainder[97]), .ZN(n4166) );
  NOR4_X2 U2290 ( .A1(remainder[93]), .A2(remainder[92]), .A3(remainder[91]), 
        .A4(remainder[90]), .ZN(n4164) );
  NOR4_X2 U2292 ( .A1(n4167), .A2(n4168), .A3(n4169), .A4(n4170), .ZN(n4145)
         );
  NAND4_X2 U2293 ( .A1(n4171), .A2(n4172), .A3(n4173), .A4(n4174), .ZN(n4170)
         );
  NOR4_X2 U2294 ( .A1(remainder[13]), .A2(remainder[12]), .A3(remainder[11]), 
        .A4(remainder[10]), .ZN(n4174) );
  NAND4_X2 U2298 ( .A1(n4175), .A2(n4176), .A3(n4177), .A4(n4178), .ZN(n4169)
         );
  NOR4_X2 U2299 ( .A1(remainder[26]), .A2(remainder[25]), .A3(remainder[24]), 
        .A4(remainder[23]), .ZN(n4178) );
  NOR4_X2 U2301 ( .A1(remainder[1]), .A2(remainder[19]), .A3(remainder[18]), 
        .A4(remainder[17]), .ZN(n4176) );
  NAND4_X2 U2303 ( .A1(n4179), .A2(n4180), .A3(n4181), .A4(n4182), .ZN(n4168)
         );
  NOR4_X2 U2304 ( .A1(remainder[38]), .A2(remainder[37]), .A3(remainder[36]), 
        .A4(remainder[35]), .ZN(n4182) );
  NAND4_X2 U2308 ( .A1(n4183), .A2(n4184), .A3(n4185), .A4(n4186), .ZN(n4167)
         );
  NOR4_X2 U2309 ( .A1(remainder[50]), .A2(remainder[4]), .A3(remainder[49]), 
        .A4(remainder[48]), .ZN(n4186) );
  NOR4_X2 U2311 ( .A1(remainder[44]), .A2(remainder[43]), .A3(remainder[42]), 
        .A4(remainder[41]), .ZN(n4184) );
  NAND2_X2 U2313 ( .A1(rmode_r3[0]), .A2(n4351), .ZN(n3741) );
  NAND2_X2 U2315 ( .A1(n2507), .A2(n4355), .ZN(n3297) );
  OAI211_X2 U2318 ( .C1(n4355), .C2(n4382), .A(n3303), .B(n4188), .ZN(n4187)
         );
  NAND2_X2 U2320 ( .A1(n4569), .A2(n4291), .ZN(n2507) );
  NAND2_X2 U2321 ( .A1(fpu_op_r3[1]), .A2(n4274), .ZN(n3973) );
  NAND2_X2 U2325 ( .A1(n2434), .A2(n4355), .ZN(n2439) );
  NAND2_X2 U2329 ( .A1(fpu_op_r3[1]), .A2(fpu_op_r3[0]), .ZN(n3458) );
  XOR2_X2 U2330 ( .A(n3065), .B(n4190), .Z(N789) );
  NAND2_X2 U2331 ( .A1(rmode_r2[1]), .A2(rmode_r2[0]), .ZN(n3065) );
  OAI221_X2 U2332 ( .B1(n4561), .B2(n4336), .C1(n4559), .C2(n5958), .A(n4554), 
        .ZN(N769) );
  OAI221_X2 U2333 ( .B1(n4561), .B2(n4335), .C1(n4560), .C2(n5959), .A(n4554), 
        .ZN(N768) );
  OAI221_X2 U2334 ( .B1(n4191), .B2(n4334), .C1(n4559), .C2(n5960), .A(n4554), 
        .ZN(N767) );
  OAI221_X2 U2335 ( .B1(n4191), .B2(n4332), .C1(n4560), .C2(n5961), .A(n4554), 
        .ZN(N766) );
  OAI221_X2 U2336 ( .B1(n4191), .B2(n4331), .C1(n4560), .C2(n5962), .A(n4554), 
        .ZN(N765) );
  OAI221_X2 U2337 ( .B1(n4191), .B2(n4333), .C1(n4560), .C2(n5963), .A(n4554), 
        .ZN(N764) );
  OAI221_X2 U2338 ( .B1(n4191), .B2(n4329), .C1(n4560), .C2(n5964), .A(n4554), 
        .ZN(N763) );
  OAI221_X2 U2339 ( .B1(n4191), .B2(n4483), .C1(n4560), .C2(n5965), .A(n4554), 
        .ZN(N762) );
  OAI221_X2 U2340 ( .B1(n4191), .B2(n4532), .C1(n4560), .C2(n5966), .A(n4554), 
        .ZN(N761) );
  OAI221_X2 U2341 ( .B1(n4191), .B2(n4531), .C1(n4560), .C2(n5967), .A(n4554), 
        .ZN(N760) );
  OAI221_X2 U2342 ( .B1(n4561), .B2(n4530), .C1(n4560), .C2(n5968), .A(n4554), 
        .ZN(N759) );
  OAI221_X2 U2343 ( .B1(n4561), .B2(n4529), .C1(n4560), .C2(n5969), .A(n4555), 
        .ZN(N758) );
  OAI221_X2 U2344 ( .B1(n4561), .B2(n4528), .C1(n4560), .C2(n5970), .A(n4555), 
        .ZN(N757) );
  OAI221_X2 U2345 ( .B1(n4561), .B2(n4527), .C1(n4560), .C2(n5971), .A(n4555), 
        .ZN(N756) );
  OAI221_X2 U2346 ( .B1(n4561), .B2(n4526), .C1(n4559), .C2(n5972), .A(n4555), 
        .ZN(N755) );
  OAI221_X2 U2347 ( .B1(n4561), .B2(n4525), .C1(n4559), .C2(n5973), .A(n4555), 
        .ZN(N754) );
  OAI221_X2 U2348 ( .B1(n4561), .B2(n4524), .C1(n4559), .C2(n5974), .A(n4555), 
        .ZN(N753) );
  OAI221_X2 U2349 ( .B1(n4561), .B2(n4523), .C1(n4559), .C2(n5975), .A(n4555), 
        .ZN(N752) );
  OAI221_X2 U2350 ( .B1(n4561), .B2(n4522), .C1(n4559), .C2(n5976), .A(n4555), 
        .ZN(N751) );
  OAI221_X2 U2351 ( .B1(n4561), .B2(n4521), .C1(n4559), .C2(n5977), .A(n4555), 
        .ZN(N750) );
  OAI221_X2 U2352 ( .B1(n4561), .B2(n4520), .C1(n4559), .C2(n5978), .A(n4555), 
        .ZN(N749) );
  OAI221_X2 U2353 ( .B1(n4561), .B2(n4519), .C1(n4559), .C2(n5979), .A(n4555), 
        .ZN(N748) );
  OAI221_X2 U2354 ( .B1(n4561), .B2(n4518), .C1(n4559), .C2(n5980), .A(n4556), 
        .ZN(N747) );
  OAI221_X2 U2355 ( .B1(n4561), .B2(n4517), .C1(n4559), .C2(n5981), .A(n4556), 
        .ZN(N746) );
  OAI221_X2 U2356 ( .B1(n4561), .B2(n4516), .C1(n4559), .C2(n5982), .A(n4556), 
        .ZN(N745) );
  OAI221_X2 U2357 ( .B1(n4561), .B2(n4515), .C1(n4558), .C2(n5983), .A(n4556), 
        .ZN(N744) );
  OAI221_X2 U2358 ( .B1(n4561), .B2(n4514), .C1(n4557), .C2(n5984), .A(n4556), 
        .ZN(N743) );
  OAI221_X2 U2359 ( .B1(n4561), .B2(n4513), .C1(n4558), .C2(n5985), .A(n4556), 
        .ZN(N742) );
  OAI221_X2 U2360 ( .B1(n4561), .B2(n4512), .C1(n4557), .C2(n5986), .A(n4556), 
        .ZN(N741) );
  OAI221_X2 U2361 ( .B1(n4561), .B2(n4511), .C1(n4558), .C2(n5987), .A(n4556), 
        .ZN(N740) );
  OAI221_X2 U2362 ( .B1(n4561), .B2(n4510), .C1(n4557), .C2(n5988), .A(n4556), 
        .ZN(N739) );
  OAI221_X2 U2363 ( .B1(n4561), .B2(n4509), .C1(n4558), .C2(n5989), .A(n4556), 
        .ZN(N738) );
  OAI221_X2 U2364 ( .B1(n4561), .B2(n4508), .C1(n4557), .C2(n5990), .A(n4556), 
        .ZN(N737) );
  OAI221_X2 U2365 ( .B1(n4561), .B2(n4507), .C1(n4558), .C2(n5991), .A(n4554), 
        .ZN(N736) );
  OAI221_X2 U2366 ( .B1(n4561), .B2(n4506), .C1(n4557), .C2(n5992), .A(n4555), 
        .ZN(N735) );
  OAI221_X2 U2367 ( .B1(n4561), .B2(n4505), .C1(n4558), .C2(n5993), .A(n4556), 
        .ZN(N734) );
  OAI221_X2 U2368 ( .B1(n4561), .B2(n4504), .C1(n4558), .C2(n5994), .A(n4554), 
        .ZN(N733) );
  OAI221_X2 U2369 ( .B1(n4561), .B2(n4503), .C1(n4558), .C2(n5995), .A(n4555), 
        .ZN(N732) );
  OAI221_X2 U2370 ( .B1(n4561), .B2(n4502), .C1(n4558), .C2(n5996), .A(n4556), 
        .ZN(N731) );
  OAI221_X2 U2371 ( .B1(n4561), .B2(n4501), .C1(n4558), .C2(n5997), .A(n4554), 
        .ZN(N730) );
  OAI221_X2 U2372 ( .B1(n4561), .B2(n4500), .C1(n4558), .C2(n5998), .A(n4555), 
        .ZN(N729) );
  OAI221_X2 U2373 ( .B1(n4561), .B2(n4499), .C1(n4558), .C2(n5999), .A(n4556), 
        .ZN(N728) );
  OAI221_X2 U2374 ( .B1(n4561), .B2(n4498), .C1(n4558), .C2(n6000), .A(n4554), 
        .ZN(N727) );
  OAI221_X2 U2375 ( .B1(n4561), .B2(n4497), .C1(n4558), .C2(n6001), .A(n4555), 
        .ZN(N726) );
  OAI221_X2 U2376 ( .B1(n4191), .B2(n4397), .C1(n4558), .C2(n6002), .A(n4556), 
        .ZN(N725) );
  OAI221_X2 U2377 ( .B1(n4191), .B2(n4396), .C1(n4558), .C2(n6003), .A(n4554), 
        .ZN(N724) );
  OAI221_X2 U2378 ( .B1(n4191), .B2(n4395), .C1(n4558), .C2(n6004), .A(n4555), 
        .ZN(N723) );
  OAI221_X2 U2379 ( .B1(n4191), .B2(n4394), .C1(n4557), .C2(n6005), .A(n4554), 
        .ZN(N722) );
  OAI221_X2 U2380 ( .B1(n4191), .B2(n4393), .C1(n4557), .C2(n6006), .A(n4556), 
        .ZN(N721) );
  OAI221_X2 U2381 ( .B1(n4191), .B2(n4392), .C1(n4557), .C2(n6007), .A(n4554), 
        .ZN(N720) );
  OAI221_X2 U2382 ( .B1(n4191), .B2(n4391), .C1(n4557), .C2(n6008), .A(n4555), 
        .ZN(N719) );
  OAI221_X2 U2383 ( .B1(n4191), .B2(n4390), .C1(n4557), .C2(n6009), .A(n4555), 
        .ZN(N718) );
  OAI221_X2 U2384 ( .B1(n4191), .B2(n4389), .C1(n4557), .C2(n6010), .A(n4556), 
        .ZN(N717) );
  OAI221_X2 U2386 ( .B1(n4191), .B2(n4388), .C1(n4557), .C2(n6011), .A(n4195), 
        .ZN(N716) );
  AOI22_X2 U2387 ( .A1(n4552), .A2(N340), .B1(N395), .B2(n4197), .ZN(n4195) );
  OAI221_X2 U2388 ( .B1(n4191), .B2(n4387), .C1(n4557), .C2(n6012), .A(n4198), 
        .ZN(N715) );
  AOI22_X2 U2389 ( .A1(n4552), .A2(opa_r1[51]), .B1(N394), .B2(n4197), .ZN(
        n4198) );
  OAI221_X2 U2390 ( .B1(n4191), .B2(n4386), .C1(n4557), .C2(n6013), .A(n4199), 
        .ZN(N714) );
  AOI22_X2 U2391 ( .A1(n4551), .A2(opa_r1[50]), .B1(N393), .B2(n4197), .ZN(
        n4199) );
  OAI221_X2 U2392 ( .B1(n4191), .B2(n4385), .C1(n4557), .C2(n6014), .A(n4200), 
        .ZN(N713) );
  AOI22_X2 U2393 ( .A1(n4552), .A2(opa_r1[49]), .B1(N392), .B2(n4197), .ZN(
        n4200) );
  OAI221_X2 U2394 ( .B1(n4191), .B2(n4496), .C1(n4557), .C2(n4380), .A(n4201), 
        .ZN(N712) );
  AOI22_X2 U2395 ( .A1(n4550), .A2(opa_r1[48]), .B1(N391), .B2(n4197), .ZN(
        n4201) );
  AOI22_X2 U2397 ( .A1(n4552), .A2(opa_r1[47]), .B1(N390), .B2(n4197), .ZN(
        n4202) );
  AOI22_X2 U2399 ( .A1(n4552), .A2(opa_r1[46]), .B1(N389), .B2(n4197), .ZN(
        n4203) );
  NAND2_X2 U2400 ( .A1(n4190), .A2(n6312), .ZN(n4191) );
  AOI22_X2 U2450 ( .A1(sign_fasu), .A2(n4303), .B1(sign_mul), .B2(fpu_op_r2[1]), .ZN(n4190) );
  NAND4_X2 U2451 ( .A1(n4483), .A2(n4329), .A3(n4250), .A4(n4251), .ZN(N340)
         );
  NOR4_X2 U2452 ( .A1(n4252), .A2(opa_r1[57]), .A3(opa_r1[59]), .A4(opa_r1[58]), .ZN(n4251) );
  OAI221_X2 U2455 ( .B1(n6312), .B2(n4381), .C1(n4330), .C2(n3296), .A(n4253), 
        .ZN(N337) );
  NAND2_X2 U2456 ( .A1(exp_fasu[10]), .A2(n4254), .ZN(n4253) );
  OAI221_X2 U2457 ( .B1(n6312), .B2(n4484), .C1(n4384), .C2(n3296), .A(n4255), 
        .ZN(N336) );
  NAND2_X2 U2458 ( .A1(exp_fasu[9]), .A2(n4254), .ZN(n4255) );
  OAI221_X2 U2459 ( .B1(n6312), .B2(n4328), .C1(n4489), .C2(n3296), .A(n4256), 
        .ZN(N335) );
  NAND2_X2 U2460 ( .A1(exp_fasu[8]), .A2(n4254), .ZN(n4256) );
  OAI221_X2 U2461 ( .B1(n6312), .B2(n4336), .C1(n4534), .C2(n3296), .A(n4257), 
        .ZN(N334) );
  NAND2_X2 U2462 ( .A1(exp_fasu[7]), .A2(n4254), .ZN(n4257) );
  OAI221_X2 U2463 ( .B1(n6312), .B2(n4335), .C1(n4536), .C2(n3296), .A(n4258), 
        .ZN(N333) );
  NAND2_X2 U2464 ( .A1(exp_fasu[6]), .A2(n4254), .ZN(n4258) );
  OAI221_X2 U2465 ( .B1(n6312), .B2(n4334), .C1(n4535), .C2(n3296), .A(n4259), 
        .ZN(N332) );
  NAND2_X2 U2466 ( .A1(exp_fasu[5]), .A2(n4254), .ZN(n4259) );
  OAI221_X2 U2467 ( .B1(n6312), .B2(n4332), .C1(n4537), .C2(n3296), .A(n4260), 
        .ZN(N331) );
  NAND2_X2 U2468 ( .A1(exp_fasu[4]), .A2(n4254), .ZN(n4260) );
  OAI221_X2 U2469 ( .B1(n6312), .B2(n4331), .C1(n4538), .C2(n3296), .A(n4261), 
        .ZN(N330) );
  NAND2_X2 U2470 ( .A1(exp_fasu[3]), .A2(n4254), .ZN(n4261) );
  OAI221_X2 U2473 ( .B1(n4262), .B2(n4333), .C1(n4539), .C2(n4303), .A(n4263), 
        .ZN(N329) );
  NAND2_X2 U2474 ( .A1(exp_fasu[2]), .A2(n4254), .ZN(n4263) );
  OAI221_X2 U2475 ( .B1(n4262), .B2(n4329), .C1(n4487), .C2(n4303), .A(n4264), 
        .ZN(N328) );
  NAND2_X2 U2476 ( .A1(exp_fasu[1]), .A2(n4254), .ZN(n4264) );
  OAI221_X2 U2477 ( .B1(n4262), .B2(n4483), .C1(n4383), .C2(n4303), .A(n4265), 
        .ZN(N327) );
  NAND2_X2 U2478 ( .A1(exp_fasu[0]), .A2(n4254), .ZN(n4265) );
  NAND2_X2 U2480 ( .A1(fpu_op_r2[2]), .A2(fpu_op_r2[0]), .ZN(n4262) );
  OAI33_X1 U3364 ( .A1(n6464), .A2(n2506), .A3(n2507), .B1(n2508), .B2(n2509), 
        .B3(n2510), .ZN(n2505) );
  OAI33_X1 U3366 ( .A1(n2598), .A2(n6355), .A3(n6357), .B1(n2671), .B2(n6376), 
        .B3(n6378), .ZN(n2652) );
  OAI33_X1 U3367 ( .A1(n2642), .A2(fract_denorm[81]), .A3(n6384), .B1(n6335), 
        .B2(fract_denorm[73]), .B3(n6397), .ZN(n2678) );
  OAI33_X1 U3368 ( .A1(n6334), .A2(fract_denorm[65]), .A3(n6390), .B1(n6326), 
        .B2(fract_denorm[57]), .B3(n6371), .ZN(n2677) );
  OAI33_X1 U3369 ( .A1(n2632), .A2(n6438), .A3(n2680), .B1(n6332), .B2(n6431), 
        .B3(n2681), .ZN(n2676) );
  OAI33_X1 U3370 ( .A1(n2598), .A2(fract_denorm[97]), .A3(n6356), .B1(n2671), 
        .B2(fract_denorm[89]), .B3(n6377), .ZN(n2687) );
  OAI33_X1 U3371 ( .A1(n3090), .A2(fracta_mul[2]), .A3(fracta_mul[1]), .B1(
        n3248), .B2(fracta_mul[17]), .B3(n4362), .ZN(n3247) );
  OAI33_X1 U3372 ( .A1(n6295), .A2(fracta_mul[47]), .A3(n4477), .B1(n6293), 
        .B2(fracta_mul[43]), .B3(n4286), .ZN(n3250) );
  OAI33_X1 U3373 ( .A1(n4372), .A2(fracta_mul[15]), .A3(n6300), .B1(n4300), 
        .B2(fracta_mul[11]), .B3(n6302), .ZN(n3274) );
  OAI33_X1 U3374 ( .A1(n6293), .A2(n6297), .A3(n4478), .B1(n3284), .B2(n3288), 
        .B3(n4376), .ZN(n3227) );
  OAI33_X1 U3375 ( .A1(n6449), .A2(n3342), .A3(n4274), .B1(n3343), .B2(
        inf_mul_r), .B3(n3344), .ZN(N902) );
  OAI33_X1 U3376 ( .A1(n3343), .A2(inf_d), .A3(n3454), .B1(n3455), .B2(
        fpu_op_r3[2]), .B3(n3456), .ZN(N899) );
  OAI33_X1 U3377 ( .A1(n3473), .A2(n2422), .A3(n4452), .B1(n3474), .B2(n6466), 
        .B3(n3475), .ZN(n3472) );
  OAI33_X1 U3378 ( .A1(n3783), .A2(u4_N6410), .A3(n4355), .B1(n4351), .B2(sign), .B3(n3784), .ZN(n3478) );
  DFF_X2 opa_r_reg_63_ ( .D(opa[63]), .CK(clk), .Q(opa_r[63]), .QN(n4533) );
  DFF_X2 opa_r_reg_62_ ( .D(opa[62]), .CK(clk), .Q(opa_r[62]), .QN(n4458) );
  DFF_X2 opa_r_reg_61_ ( .D(opa[61]), .CK(clk), .Q(opa_r[61]), .QN(n4448) );
  DFF_X2 opa_r_reg_60_ ( .D(opa[60]), .CK(clk), .Q(opa_r[60]), .QN(n4357) );
  DFF_X2 opa_r_reg_59_ ( .D(opa[59]), .CK(clk), .Q(opa_r[59]), .QN(n4442) );
  DFF_X2 opa_r_reg_58_ ( .D(opa[58]), .CK(clk), .Q(opa_r[58]), .QN(n4454) );
  DFF_X2 opa_r_reg_57_ ( .D(opa[57]), .CK(clk), .Q(opa_r[57]), .QN(n4453) );
  DFF_X2 opa_r_reg_56_ ( .D(opa[56]), .CK(clk), .Q(opa_r[56]), .QN(n4456) );
  DFF_X2 opa_r_reg_55_ ( .D(opa[55]), .CK(clk), .Q(opa_r[55]), .QN(n4358) );
  DFF_X2 opa_r_reg_54_ ( .D(opa[54]), .CK(clk), .Q(opa_r[54]), .QN(n4451) );
  DFF_X2 opa_r_reg_53_ ( .D(opa[53]), .CK(clk), .Q(opa_r[53]), .QN(n4450) );
  DFF_X2 opa_r_reg_52_ ( .D(opa[52]), .CK(clk), .Q(opa_r[52]), .QN(n4449) );
  DFF_X2 opa_r_reg_51_ ( .D(opa[51]), .CK(clk), .Q(fracta_mul[51]), .QN(n4273)
         );
  DFF_X2 opa_r_reg_50_ ( .D(opa[50]), .CK(clk), .Q(fracta_mul[50]), .QN(n4480)
         );
  DFF_X2 opa_r_reg_49_ ( .D(opa[49]), .CK(clk), .Q(fracta_mul[49]) );
  DFF_X2 opa_r_reg_48_ ( .D(opa[48]), .CK(clk), .Q(fracta_mul[48]) );
  DFF_X2 opa_r_reg_47_ ( .D(opa[47]), .CK(clk), .Q(fracta_mul[47]) );
  DFF_X2 opa_r_reg_46_ ( .D(opa[46]), .CK(clk), .Q(fracta_mul[46]), .QN(n4477)
         );
  DFF_X2 opa_r_reg_45_ ( .D(opa[45]), .CK(clk), .Q(fracta_mul[45]), .QN(n4367)
         );
  DFF_X2 opa_r_reg_44_ ( .D(opa[44]), .CK(clk), .Q(fracta_mul[44]), .QN(n4277)
         );
  DFF_X2 opa_r_reg_43_ ( .D(opa[43]), .CK(clk), .Q(fracta_mul[43]) );
  DFF_X2 opa_r_reg_42_ ( .D(opa[42]), .CK(clk), .Q(fracta_mul[42]), .QN(n4286)
         );
  DFF_X2 opa_r_reg_41_ ( .D(opa[41]), .CK(clk), .Q(fracta_mul[41]), .QN(n4472)
         );
  DFF_X2 opa_r_reg_40_ ( .D(opa[40]), .CK(clk), .Q(fracta_mul[40]) );
  DFF_X2 opa_r_reg_39_ ( .D(opa[39]), .CK(clk), .Q(fracta_mul[39]), .QN(n4478)
         );
  DFF_X2 opa_r_reg_38_ ( .D(opa[38]), .CK(clk), .Q(fracta_mul[38]), .QN(n4284)
         );
  DFF_X2 opa_r_reg_37_ ( .D(opa[37]), .CK(clk), .Q(fracta_mul[37]), .QN(n4272)
         );
  DFF_X2 opa_r_reg_36_ ( .D(opa[36]), .CK(clk), .Q(fracta_mul[36]), .QN(n4276)
         );
  DFF_X2 opa_r_reg_35_ ( .D(opa[35]), .CK(clk), .Q(fracta_mul[35]), .QN(n4474)
         );
  DFF_X2 opa_r_reg_34_ ( .D(opa[34]), .CK(clk), .Q(fracta_mul[34]) );
  DFF_X2 opa_r_reg_33_ ( .D(opa[33]), .CK(clk), .Q(fracta_mul[33]) );
  DFF_X2 opa_r_reg_32_ ( .D(opa[32]), .CK(clk), .Q(fracta_mul[32]), .QN(n4287)
         );
  DFF_X2 opa_r_reg_31_ ( .D(opa[31]), .CK(clk), .Q(fracta_mul[31]), .QN(n4370)
         );
  DFF_X2 opa_r_reg_30_ ( .D(opa[30]), .CK(clk), .Q(fracta_mul[30]), .QN(n4479)
         );
  DFF_X2 opa_r_reg_29_ ( .D(opa[29]), .CK(clk), .Q(fracta_mul[29]), .QN(n4475)
         );
  DFF_X2 opa_r_reg_28_ ( .D(opa[28]), .CK(clk), .Q(fracta_mul[28]), .QN(n4285)
         );
  DFF_X2 opa_r_reg_27_ ( .D(opa[27]), .CK(clk), .Q(fracta_mul[27]), .QN(n4301)
         );
  DFF_X2 opa_r_reg_26_ ( .D(opa[26]), .CK(clk), .Q(fracta_mul[26]) );
  DFF_X2 opa_r_reg_25_ ( .D(opa[25]), .CK(clk), .Q(fracta_mul[25]), .QN(n4473)
         );
  DFF_X2 opa_r_reg_24_ ( .D(opa[24]), .CK(clk), .Q(fracta_mul[24]) );
  DFF_X2 opa_r_reg_23_ ( .D(opa[23]), .CK(clk), .Q(fracta_mul[23]) );
  DFF_X2 opa_r_reg_22_ ( .D(opa[22]), .CK(clk), .Q(fracta_mul[22]), .QN(n4283)
         );
  DFF_X2 opa_r_reg_21_ ( .D(opa[21]), .CK(clk), .Q(fracta_mul[21]), .QN(n4292)
         );
  DFF_X2 opa_r_reg_20_ ( .D(opa[20]), .CK(clk), .Q(fracta_mul[20]), .QN(n4320)
         );
  DFF_X2 opa_r_reg_19_ ( .D(opa[19]), .CK(clk), .Q(fracta_mul[19]) );
  DFF_X2 opa_r_reg_18_ ( .D(opa[18]), .CK(clk), .Q(fracta_mul[18]), .QN(n4369)
         );
  DFF_X2 opa_r_reg_17_ ( .D(opa[17]), .CK(clk), .Q(fracta_mul[17]), .QN(n4319)
         );
  DFF_X2 opa_r_reg_16_ ( .D(opa[16]), .CK(clk), .Q(fracta_mul[16]), .QN(n4362)
         );
  DFF_X2 opa_r_reg_15_ ( .D(opa[15]), .CK(clk), .Q(fracta_mul[15]), .QN(n4318)
         );
  DFF_X2 opa_r_reg_14_ ( .D(opa[14]), .CK(clk), .Q(fracta_mul[14]), .QN(n4372)
         );
  DFF_X2 opa_r_reg_13_ ( .D(opa[13]), .CK(clk), .Q(fracta_mul[13]), .QN(n4476)
         );
  DFF_X2 opa_r_reg_12_ ( .D(opa[12]), .CK(clk), .Q(fracta_mul[12]), .QN(n4374)
         );
  DFF_X2 opa_r_reg_11_ ( .D(opa[11]), .CK(clk), .Q(fracta_mul[11]), .QN(n4361)
         );
  DFF_X2 opa_r_reg_10_ ( .D(opa[10]), .CK(clk), .Q(fracta_mul[10]), .QN(n4300)
         );
  DFF_X2 opa_r_reg_9_ ( .D(opa[9]), .CK(clk), .Q(fracta_mul[9]), .QN(n4368) );
  DFF_X2 opa_r_reg_8_ ( .D(opa[8]), .CK(clk), .Q(fracta_mul[8]), .QN(n4326) );
  DFF_X2 opa_r_reg_7_ ( .D(opa[7]), .CK(clk), .Q(fracta_mul[7]), .QN(n4376) );
  DFF_X2 opa_r_reg_6_ ( .D(opa[6]), .CK(clk), .Q(fracta_mul[6]), .QN(n4375) );
  DFF_X2 opa_r_reg_5_ ( .D(opa[5]), .CK(clk), .Q(fracta_mul[5]), .QN(n4371) );
  DFF_X2 opa_r_reg_4_ ( .D(opa[4]), .CK(clk), .Q(fracta_mul[4]) );
  DFF_X2 opa_r_reg_3_ ( .D(opa[3]), .CK(clk), .Q(fracta_mul[3]), .QN(n4360) );
  DFF_X2 opa_r_reg_2_ ( .D(opa[2]), .CK(clk), .Q(fracta_mul[2]) );
  DFF_X2 opa_r_reg_1_ ( .D(opa[1]), .CK(clk), .Q(fracta_mul[1]), .QN(n4373) );
  DFF_X2 opa_r_reg_0_ ( .D(opa[0]), .CK(clk), .Q(fracta_mul[0]), .QN(n4322) );
  DFF_X2 opb_r_reg_63_ ( .D(opb[63]), .CK(clk), .Q(opb_r[63]) );
  DFF_X2 opb_r_reg_62_ ( .D(opb[62]), .CK(clk), .Q(opb_r[62]), .QN(n4363) );
  DFF_X2 opb_r_reg_61_ ( .D(opb[61]), .CK(clk), .Q(opb_r[61]) );
  DFF_X2 opb_r_reg_60_ ( .D(opb[60]), .CK(clk), .Q(opb_r[60]) );
  DFF_X2 opb_r_reg_59_ ( .D(opb[59]), .CK(clk), .Q(opb_r[59]), .QN(n4340) );
  DFF_X2 opb_r_reg_58_ ( .D(opb[58]), .CK(clk), .Q(opb_r[58]), .QN(n4399) );
  DFF_X2 opb_r_reg_57_ ( .D(opb[57]), .CK(clk), .Q(opb_r[57]), .QN(n4296) );
  DFF_X2 opb_r_reg_56_ ( .D(opb[56]), .CK(clk), .Q(opb_r[56]), .QN(n4359) );
  DFF_X2 opb_r_reg_55_ ( .D(opb[55]), .CK(clk), .Q(opb_r[55]), .QN(n4321) );
  DFF_X2 opb_r_reg_54_ ( .D(opb[54]), .CK(clk), .Q(opb_r[54]), .QN(n4457) );
  DFF_X2 opb_r_reg_53_ ( .D(opb[53]), .CK(clk), .Q(opb_r[53]), .QN(n4275) );
  DFF_X2 opb_r_reg_52_ ( .D(opb[52]), .CK(clk), .Q(opb_r[52]), .QN(n4270) );
  DFF_X2 opb_r_reg_51_ ( .D(opb[51]), .CK(clk), .Q(u6_N51), .QN(n4459) );
  DFF_X2 opb_r_reg_50_ ( .D(opb[50]), .CK(clk), .Q(u6_N50) );
  DFF_X2 opb_r_reg_49_ ( .D(opb[49]), .CK(clk), .Q(u6_N49) );
  DFF_X2 opb_r_reg_48_ ( .D(opb[48]), .CK(clk), .Q(u6_N48) );
  DFF_X2 opb_r_reg_47_ ( .D(opb[47]), .CK(clk), .Q(u6_N47) );
  DFF_X2 opb_r_reg_46_ ( .D(opb[46]), .CK(clk), .Q(u6_N46) );
  DFF_X2 opb_r_reg_45_ ( .D(opb[45]), .CK(clk), .Q(u6_N45) );
  DFF_X2 opb_r_reg_44_ ( .D(opb[44]), .CK(clk), .Q(u6_N44), .QN(n4468) );
  DFF_X2 opb_r_reg_43_ ( .D(opb[43]), .CK(clk), .Q(u6_N43) );
  DFF_X2 opb_r_reg_42_ ( .D(opb[42]), .CK(clk), .Q(u6_N42), .QN(n4467) );
  DFF_X2 opb_r_reg_41_ ( .D(opb[41]), .CK(clk), .Q(u6_N41) );
  DFF_X2 opb_r_reg_40_ ( .D(opb[40]), .CK(clk), .Q(u6_N40) );
  DFF_X2 opb_r_reg_39_ ( .D(opb[39]), .CK(clk), .Q(u6_N39) );
  DFF_X2 opb_r_reg_38_ ( .D(opb[38]), .CK(clk), .Q(u6_N38), .QN(n4465) );
  DFF_X2 opb_r_reg_37_ ( .D(opb[37]), .CK(clk), .Q(u6_N37), .QN(n4471) );
  DFF_X2 opb_r_reg_36_ ( .D(opb[36]), .CK(clk), .Q(u6_N36), .QN(n4470) );
  DFF_X2 opb_r_reg_35_ ( .D(opb[35]), .CK(clk), .Q(u6_N35) );
  DFF_X2 opb_r_reg_34_ ( .D(opb[34]), .CK(clk), .Q(u6_N34) );
  DFF_X2 opb_r_reg_33_ ( .D(opb[33]), .CK(clk), .Q(u6_N33) );
  DFF_X2 opb_r_reg_32_ ( .D(opb[32]), .CK(clk), .Q(u6_N32), .QN(n4464) );
  DFF_X2 opb_r_reg_31_ ( .D(opb[31]), .CK(clk), .Q(u6_N31) );
  DFF_X2 opb_r_reg_30_ ( .D(opb[30]), .CK(clk), .Q(u6_N30) );
  DFF_X2 opb_r_reg_29_ ( .D(opb[29]), .CK(clk), .Q(u6_N29) );
  DFF_X2 opb_r_reg_28_ ( .D(opb[28]), .CK(clk), .Q(u6_N28), .QN(n4469) );
  DFF_X2 opb_r_reg_27_ ( .D(opb[27]), .CK(clk), .Q(u6_N27), .QN(n4466) );
  DFF_X2 opb_r_reg_26_ ( .D(opb[26]), .CK(clk), .Q(u6_N26) );
  DFF_X2 opb_r_reg_25_ ( .D(opb[25]), .CK(clk), .Q(u6_N25) );
  DFF_X2 opb_r_reg_24_ ( .D(opb[24]), .CK(clk), .Q(u6_N24) );
  DFF_X2 opb_r_reg_23_ ( .D(opb[23]), .CK(clk), .Q(u6_N23) );
  DFF_X2 opb_r_reg_22_ ( .D(opb[22]), .CK(clk), .Q(u6_N22), .QN(n4462) );
  DFF_X2 opb_r_reg_21_ ( .D(opb[21]), .CK(clk), .Q(u6_N21), .QN(n4325) );
  DFF_X2 opb_r_reg_20_ ( .D(opb[20]), .CK(clk), .Q(u6_N20), .QN(n4366) );
  DFF_X2 opb_r_reg_19_ ( .D(opb[19]), .CK(clk), .Q(u6_N19) );
  DFF_X2 opb_r_reg_18_ ( .D(opb[18]), .CK(clk), .Q(u6_N18) );
  DFF_X2 opb_r_reg_17_ ( .D(opb[17]), .CK(clk), .Q(u6_N17), .QN(n4461) );
  DFF_X2 opb_r_reg_16_ ( .D(opb[16]), .CK(clk), .Q(u6_N16), .QN(n4324) );
  DFF_X2 opb_r_reg_15_ ( .D(opb[15]), .CK(clk), .Q(u6_N15), .QN(n4365) );
  DFF_X2 opb_r_reg_14_ ( .D(opb[14]), .CK(clk), .Q(u6_N14) );
  DFF_X2 opb_r_reg_13_ ( .D(opb[13]), .CK(clk), .Q(u6_N13) );
  DFF_X2 opb_r_reg_12_ ( .D(opb[12]), .CK(clk), .Q(u6_N12) );
  DFF_X2 opb_r_reg_11_ ( .D(opb[11]), .CK(clk), .Q(u6_N11), .QN(n4460) );
  DFF_X2 opb_r_reg_10_ ( .D(opb[10]), .CK(clk), .Q(u6_N10), .QN(n4323) );
  DFF_X2 opb_r_reg_9_ ( .D(opb[9]), .CK(clk), .Q(u6_N9) );
  DFF_X2 opb_r_reg_8_ ( .D(opb[8]), .CK(clk), .Q(u6_N8) );
  DFF_X2 opb_r_reg_7_ ( .D(opb[7]), .CK(clk), .Q(u6_N7) );
  DFF_X2 opb_r_reg_6_ ( .D(opb[6]), .CK(clk), .Q(u6_N6) );
  DFF_X2 opb_r_reg_5_ ( .D(opb[5]), .CK(clk), .Q(u6_N5) );
  DFF_X2 opb_r_reg_4_ ( .D(opb[4]), .CK(clk), .Q(u6_N4) );
  DFF_X2 opb_r_reg_3_ ( .D(opb[3]), .CK(clk), .Q(u6_N3), .QN(n4463) );
  DFF_X2 opb_r_reg_2_ ( .D(opb[2]), .CK(clk), .Q(u6_N2) );
  DFF_X2 opb_r_reg_1_ ( .D(opb[1]), .CK(clk), .Q(u6_N1) );
  DFF_X2 opb_r_reg_0_ ( .D(opb[0]), .CK(clk), .Q(u6_N0), .QN(n4364) );
  DFF_X2 rmode_r1_reg_1_ ( .D(rmode[1]), .CK(clk), .Q(rmode_r1[1]) );
  DFF_X2 rmode_r1_reg_0_ ( .D(rmode[0]), .CK(clk), .Q(rmode_r1[0]) );
  DFF_X2 rmode_r2_reg_1_ ( .D(rmode_r1[1]), .CK(clk), .Q(rmode_r2[1]) );
  DFF_X2 rmode_r2_reg_0_ ( .D(rmode_r1[0]), .CK(clk), .Q(rmode_r2[0]) );
  DFF_X2 rmode_r3_reg_1_ ( .D(rmode_r2[1]), .CK(clk), .Q(rmode_r3[1]), .QN(
        n4351) );
  DFF_X2 rmode_r3_reg_0_ ( .D(rmode_r2[0]), .CK(clk), .Q(rmode_r3[0]), .QN(
        n4441) );
  DFF_X2 fpu_op_r1_reg_2_ ( .D(fpu_op[2]), .CK(clk), .Q(fpu_op_r1[2]), .QN(
        n4377) );
  DFF_X2 fpu_op_r1_reg_1_ ( .D(fpu_op[1]), .CK(clk), .Q(fpu_op_r1[1]) );
  DFF_X2 fpu_op_r1_reg_0_ ( .D(fpu_op[0]), .CK(clk), .Q(fpu_op_r1[0]), .QN(
        n4481) );
  DFF_X2 fpu_op_r2_reg_2_ ( .D(fpu_op_r1[2]), .CK(clk), .Q(fpu_op_r2[2]) );
  DFF_X2 fpu_op_r2_reg_1_ ( .D(fpu_op_r1[1]), .CK(clk), .Q(fpu_op_r2[1]), .QN(
        n4303) );
  DFF_X2 fpu_op_r2_reg_0_ ( .D(fpu_op_r1[0]), .CK(clk), .Q(fpu_op_r2[0]), .QN(
        n4493) );
  DFF_X2 fpu_op_r3_reg_2_ ( .D(fpu_op_r2[2]), .CK(clk), .Q(fpu_op_r3[2]), .QN(
        n4291) );
  DFF_X2 fpu_op_r3_reg_1_ ( .D(fpu_op_r2[1]), .CK(clk), .Q(fpu_op_r3[1]), .QN(
        n4400) );
  DFF_X2 fpu_op_r3_reg_0_ ( .D(fpu_op_r2[0]), .CK(clk), .Q(fpu_op_r3[0]), .QN(
        n4274) );
  DFF_X2 div_opa_ldz_r1_reg_4_ ( .D(div_opa_ldz_d[4]), .CK(clk), .Q(
        div_opa_ldz_r1[4]) );
  DFF_X2 div_opa_ldz_r1_reg_3_ ( .D(div_opa_ldz_d[3]), .CK(clk), .Q(
        div_opa_ldz_r1[3]) );
  DFF_X2 div_opa_ldz_r1_reg_2_ ( .D(div_opa_ldz_d[2]), .CK(clk), .Q(
        div_opa_ldz_r1[2]) );
  DFF_X2 div_opa_ldz_r1_reg_1_ ( .D(div_opa_ldz_d[1]), .CK(clk), .Q(
        div_opa_ldz_r1[1]) );
  DFF_X2 div_opa_ldz_r1_reg_0_ ( .D(div_opa_ldz_d[0]), .CK(clk), .Q(
        div_opa_ldz_r1[0]) );
  DFF_X2 div_opa_ldz_r2_reg_4_ ( .D(div_opa_ldz_r1[4]), .CK(clk), .Q(
        div_opa_ldz_r2[4]), .QN(n4445) );
  DFF_X2 div_opa_ldz_r2_reg_3_ ( .D(div_opa_ldz_r1[3]), .CK(clk), .Q(
        div_opa_ldz_r2[3]), .QN(n4443) );
  DFF_X2 div_opa_ldz_r2_reg_2_ ( .D(div_opa_ldz_r1[2]), .CK(clk), .Q(
        div_opa_ldz_r2[2]), .QN(n4444) );
  DFF_X2 div_opa_ldz_r2_reg_1_ ( .D(div_opa_ldz_r1[1]), .CK(clk), .Q(
        div_opa_ldz_r2[1]), .QN(n4446) );
  DFF_X2 div_opa_ldz_r2_reg_0_ ( .D(div_opa_ldz_r1[0]), .CK(clk), .Q(
        div_opa_ldz_r2[0]), .QN(n4447) );
  DFF_X2 opa_r1_reg_62_ ( .D(opa_r[62]), .CK(clk), .QN(n4381) );
  DFF_X2 opa_r1_reg_61_ ( .D(opa_r[61]), .CK(clk), .QN(n4484) );
  DFF_X2 opa_r1_reg_60_ ( .D(opa_r[60]), .CK(clk), .QN(n4328) );
  DFF_X2 opa_r1_reg_59_ ( .D(opa_r[59]), .CK(clk), .Q(opa_r1[59]), .QN(n4336)
         );
  DFF_X2 opa_r1_reg_58_ ( .D(opa_r[58]), .CK(clk), .Q(opa_r1[58]), .QN(n4335)
         );
  DFF_X2 opa_r1_reg_57_ ( .D(opa_r[57]), .CK(clk), .Q(opa_r1[57]), .QN(n4334)
         );
  DFF_X2 opa_r1_reg_56_ ( .D(opa_r[56]), .CK(clk), .Q(opa_r1[56]), .QN(n4332)
         );
  DFF_X2 opa_r1_reg_55_ ( .D(opa_r[55]), .CK(clk), .Q(opa_r1[55]), .QN(n4331)
         );
  DFF_X2 opa_r1_reg_54_ ( .D(opa_r[54]), .CK(clk), .Q(opa_r1[54]), .QN(n4333)
         );
  DFF_X2 opa_r1_reg_53_ ( .D(opa_r[53]), .CK(clk), .Q(opa_r1[53]), .QN(n4329)
         );
  DFF_X2 opa_r1_reg_52_ ( .D(opa_r[52]), .CK(clk), .Q(opa_r1[52]), .QN(n4483)
         );
  DFF_X2 opa_r1_reg_51_ ( .D(fracta_mul[51]), .CK(clk), .Q(opa_r1[51]), .QN(
        n4532) );
  DFF_X2 opa_r1_reg_50_ ( .D(fracta_mul[50]), .CK(clk), .Q(opa_r1[50]), .QN(
        n4531) );
  DFF_X2 opa_r1_reg_49_ ( .D(fracta_mul[49]), .CK(clk), .Q(opa_r1[49]), .QN(
        n4530) );
  DFF_X2 opa_r1_reg_48_ ( .D(fracta_mul[48]), .CK(clk), .Q(opa_r1[48]), .QN(
        n4529) );
  DFF_X2 opa_r1_reg_47_ ( .D(fracta_mul[47]), .CK(clk), .Q(opa_r1[47]), .QN(
        n4528) );
  DFF_X2 opa_r1_reg_46_ ( .D(fracta_mul[46]), .CK(clk), .Q(opa_r1[46]), .QN(
        n4527) );
  DFF_X2 opa_r1_reg_45_ ( .D(fracta_mul[45]), .CK(clk), .Q(opa_r1[45]), .QN(
        n4526) );
  DFF_X2 opa_r1_reg_44_ ( .D(fracta_mul[44]), .CK(clk), .Q(opa_r1[44]), .QN(
        n4525) );
  DFF_X2 opa_r1_reg_43_ ( .D(fracta_mul[43]), .CK(clk), .Q(opa_r1[43]), .QN(
        n4524) );
  DFF_X2 opa_r1_reg_42_ ( .D(fracta_mul[42]), .CK(clk), .Q(opa_r1[42]), .QN(
        n4523) );
  DFF_X2 opa_r1_reg_41_ ( .D(fracta_mul[41]), .CK(clk), .Q(opa_r1[41]), .QN(
        n4522) );
  DFF_X2 opa_r1_reg_40_ ( .D(fracta_mul[40]), .CK(clk), .Q(opa_r1[40]), .QN(
        n4521) );
  DFF_X2 opa_r1_reg_39_ ( .D(fracta_mul[39]), .CK(clk), .Q(opa_r1[39]), .QN(
        n4520) );
  DFF_X2 opa_r1_reg_38_ ( .D(fracta_mul[38]), .CK(clk), .Q(opa_r1[38]), .QN(
        n4519) );
  DFF_X2 opa_r1_reg_37_ ( .D(fracta_mul[37]), .CK(clk), .Q(opa_r1[37]), .QN(
        n4518) );
  DFF_X2 opa_r1_reg_36_ ( .D(fracta_mul[36]), .CK(clk), .Q(opa_r1[36]), .QN(
        n4517) );
  DFF_X2 opa_r1_reg_35_ ( .D(fracta_mul[35]), .CK(clk), .Q(opa_r1[35]), .QN(
        n4516) );
  DFF_X2 opa_r1_reg_34_ ( .D(fracta_mul[34]), .CK(clk), .Q(opa_r1[34]), .QN(
        n4515) );
  DFF_X2 opa_r1_reg_33_ ( .D(fracta_mul[33]), .CK(clk), .Q(opa_r1[33]), .QN(
        n4514) );
  DFF_X2 opa_r1_reg_32_ ( .D(fracta_mul[32]), .CK(clk), .Q(opa_r1[32]), .QN(
        n4513) );
  DFF_X2 opa_r1_reg_31_ ( .D(fracta_mul[31]), .CK(clk), .Q(opa_r1[31]), .QN(
        n4512) );
  DFF_X2 opa_r1_reg_30_ ( .D(fracta_mul[30]), .CK(clk), .Q(opa_r1[30]), .QN(
        n4511) );
  DFF_X2 opa_r1_reg_29_ ( .D(fracta_mul[29]), .CK(clk), .Q(opa_r1[29]), .QN(
        n4510) );
  DFF_X2 opa_r1_reg_28_ ( .D(fracta_mul[28]), .CK(clk), .Q(opa_r1[28]), .QN(
        n4509) );
  DFF_X2 opa_r1_reg_27_ ( .D(fracta_mul[27]), .CK(clk), .Q(opa_r1[27]), .QN(
        n4508) );
  DFF_X2 opa_r1_reg_26_ ( .D(fracta_mul[26]), .CK(clk), .Q(opa_r1[26]), .QN(
        n4507) );
  DFF_X2 opa_r1_reg_25_ ( .D(fracta_mul[25]), .CK(clk), .Q(opa_r1[25]), .QN(
        n4506) );
  DFF_X2 opa_r1_reg_24_ ( .D(fracta_mul[24]), .CK(clk), .Q(opa_r1[24]), .QN(
        n4505) );
  DFF_X2 opa_r1_reg_23_ ( .D(fracta_mul[23]), .CK(clk), .Q(opa_r1[23]), .QN(
        n4504) );
  DFF_X2 opa_r1_reg_22_ ( .D(fracta_mul[22]), .CK(clk), .Q(opa_r1[22]), .QN(
        n4503) );
  DFF_X2 opa_r1_reg_21_ ( .D(fracta_mul[21]), .CK(clk), .Q(opa_r1[21]), .QN(
        n4502) );
  DFF_X2 opa_r1_reg_20_ ( .D(fracta_mul[20]), .CK(clk), .Q(opa_r1[20]), .QN(
        n4501) );
  DFF_X2 opa_r1_reg_19_ ( .D(fracta_mul[19]), .CK(clk), .Q(opa_r1[19]), .QN(
        n4500) );
  DFF_X2 opa_r1_reg_18_ ( .D(fracta_mul[18]), .CK(clk), .Q(opa_r1[18]), .QN(
        n4499) );
  DFF_X2 opa_r1_reg_17_ ( .D(fracta_mul[17]), .CK(clk), .Q(opa_r1[17]), .QN(
        n4498) );
  DFF_X2 opa_r1_reg_16_ ( .D(fracta_mul[16]), .CK(clk), .Q(opa_r1[16]), .QN(
        n4497) );
  DFF_X2 opa_r1_reg_15_ ( .D(fracta_mul[15]), .CK(clk), .Q(opa_r1[15]), .QN(
        n4397) );
  DFF_X2 opa_r1_reg_14_ ( .D(fracta_mul[14]), .CK(clk), .Q(opa_r1[14]), .QN(
        n4396) );
  DFF_X2 opa_r1_reg_13_ ( .D(fracta_mul[13]), .CK(clk), .Q(opa_r1[13]), .QN(
        n4395) );
  DFF_X2 opa_r1_reg_12_ ( .D(fracta_mul[12]), .CK(clk), .Q(opa_r1[12]), .QN(
        n4394) );
  DFF_X2 opa_r1_reg_11_ ( .D(fracta_mul[11]), .CK(clk), .Q(opa_r1[11]), .QN(
        n4393) );
  DFF_X2 opa_r1_reg_10_ ( .D(fracta_mul[10]), .CK(clk), .Q(opa_r1[10]), .QN(
        n4392) );
  DFF_X2 opa_r1_reg_9_ ( .D(fracta_mul[9]), .CK(clk), .Q(opa_r1[9]), .QN(n4391) );
  DFF_X2 opa_r1_reg_8_ ( .D(fracta_mul[8]), .CK(clk), .Q(opa_r1[8]), .QN(n4390) );
  DFF_X2 opa_r1_reg_7_ ( .D(fracta_mul[7]), .CK(clk), .Q(opa_r1[7]), .QN(n4389) );
  DFF_X2 opa_r1_reg_6_ ( .D(fracta_mul[6]), .CK(clk), .Q(opa_r1[6]), .QN(n4388) );
  DFF_X2 opa_r1_reg_5_ ( .D(fracta_mul[5]), .CK(clk), .Q(opa_r1[5]), .QN(n4387) );
  DFF_X2 opa_r1_reg_4_ ( .D(fracta_mul[4]), .CK(clk), .Q(opa_r1[4]), .QN(n4386) );
  DFF_X2 opa_r1_reg_3_ ( .D(fracta_mul[3]), .CK(clk), .Q(opa_r1[3]), .QN(n4385) );
  DFF_X2 opa_r1_reg_2_ ( .D(fracta_mul[2]), .CK(clk), .Q(opa_r1[2]), .QN(n4496) );
  DFF_X2 opa_r1_reg_1_ ( .D(fracta_mul[1]), .CK(clk), .Q(opa_r1[1]), .QN(n4488) );
  DFF_X2 opa_r1_reg_0_ ( .D(fracta_mul[0]), .CK(clk), .Q(N343), .QN(n4380) );
  DFF_X2 opas_r1_reg ( .D(opa_r[63]), .CK(clk), .Q(opas_r1) );
  DFF_X2 opas_r2_reg ( .D(opas_r1), .CK(clk), .Q(opas_r2) );
  DFF_X2 u0_fractb_00_reg ( .D(n4268), .CK(clk), .Q(u0_fractb_00) );
  DFF_X2 u0_fracta_00_reg ( .D(n4267), .CK(clk), .Q(u0_fracta_00) );
  DFF_X2 u0_expb_00_reg ( .D(n6303), .CK(clk), .Q(u0_expb_00) );
  DFF_X2 u0_opb_dn_reg ( .D(u0_expb_00), .CK(clk), .Q(opb_dn), .QN(n4269) );
  DFF_X2 u0_opb_00_reg ( .D(u0_N17), .CK(clk), .Q(opb_00) );
  DFF_X2 u0_expa_00_reg ( .D(n4601), .CK(clk), .Q(u0_expa_00) );
  DFF_X2 u0_opa_dn_reg ( .D(u0_expa_00), .CK(clk), .QN(n4271) );
  DFF_X2 u0_opa_00_reg ( .D(u0_N16), .CK(clk), .Q(opa_00), .QN(n4486) );
  DFF_X2 u0_opb_nan_reg ( .D(u0_N11), .CK(clk), .Q(opb_nan), .QN(n4492) );
  DFF_X2 u0_opa_nan_reg ( .D(u0_N10), .CK(clk), .Q(opa_nan) );
  DFF_X2 opa_nan_r_reg ( .D(N912), .CK(clk), .Q(opa_nan_r) );
  DFF_X2 u0_snan_r_b_reg ( .D(u0_N5), .CK(clk), .Q(u0_snan_r_b) );
  DFF_X2 u0_qnan_r_b_reg ( .D(u6_N51), .CK(clk), .Q(u0_qnan_r_b) );
  DFF_X2 u0_snan_r_a_reg ( .D(u0_N4), .CK(clk), .Q(u0_snan_r_a) );
  DFF_X2 u0_qnan_r_a_reg ( .D(fracta_mul[51]), .CK(clk), .Q(u0_qnan_r_a) );
  DFF_X2 u0_infb_f_r_reg ( .D(n4268), .CK(clk), .Q(u0_infb_f_r) );
  DFF_X2 u0_infa_f_r_reg ( .D(n4267), .CK(clk), .Q(u0_infa_f_r) );
  DFF_X2 u0_expb_ff_reg ( .D(n6304), .CK(clk), .Q(u0_expb_ff) );
  DFF_X2 u0_opb_inf_reg ( .D(n6452), .CK(clk), .Q(opb_inf), .QN(n4327) );
  DFF_X2 u0_expa_ff_reg ( .D(n6276), .CK(clk), .Q(u0_expa_ff) );
  DFF_X2 u0_snan_reg ( .D(n6450), .CK(clk), .Q(snan_d) );
  DFF_X2 snan_reg ( .D(snan_d), .CK(clk), .Q(snan) );
  DFF_X2 u0_qnan_reg ( .D(n6451), .CK(clk), .Q(qnan_d) );
  DFF_X2 u0_opa_inf_reg ( .D(n6453), .CK(clk), .Q(opa_inf), .QN(n4382) );
  DFF_X2 div_by_zero_reg ( .D(N913), .CK(clk), .Q(div_by_zero) );
  DFF_X2 u0_inf_reg ( .D(u0_N7), .CK(clk), .Q(inf_d) );
  DFF_X2 u0_ind_reg ( .D(u0_N6), .CK(clk), .Q(ind_d) );
  DFF_X2 u1_fasu_op_reg ( .D(u1_N232), .CK(clk), .Q(fasu_op), .QN(n4305) );
  DFF_X2 fasu_op_r1_reg ( .D(n4660), .CK(clk), .Q(fasu_op_r1) );
  DFF_X2 fasu_op_r2_reg ( .D(fasu_op_r1), .CK(clk), .Q(fasu_op_r2), .QN(n4494)
         );
  DFF_X2 qnan_reg ( .D(N904), .CK(clk), .Q(qnan) );
  DFF_X2 u1_fracta_eq_fractb_reg ( .D(u1_N220), .CK(clk), .Q(
        u1_fracta_eq_fractb) );
  DFF_X2 u1_fracta_lt_fractb_reg ( .D(u1_N219), .CK(clk), .Q(
        u1_fracta_lt_fractb) );
  DFF_X2 u1_add_r_reg ( .D(n4481), .CK(clk), .Q(u1_add_r) );
  DFF_X2 u1_signb_r_reg ( .D(opb_r[63]), .CK(clk), .Q(u1_signb_r), .QN(n4495)
         );
  DFF_X2 u1_signa_r_reg ( .D(opa_r[63]), .CK(clk), .Q(u1_signa_r), .QN(n4490)
         );
  DFF_X2 u1_result_zero_sign_reg ( .D(u1_N218), .CK(clk), .Q(
        result_zero_sign_d) );
  DFF_X2 u1_nan_sign_reg ( .D(u1_N229), .CK(clk), .Q(nan_sign_d) );
  DFF_X2 u1_sign_reg ( .D(u1_sign_d), .CK(clk), .Q(sign_fasu) );
  DFF_X2 sign_fasu_r_reg ( .D(sign_fasu), .CK(clk), .Q(sign_fasu_r) );
  DFF_X2 u1_fractb_out_reg_0_ ( .D(u1_fractb_s[0]), .CK(clk), .Q(fractb[0]) );
  DFF_X2 u1_fractb_out_reg_1_ ( .D(u1_fractb_s[1]), .CK(clk), .Q(fractb[1]) );
  DFF_X2 u1_fractb_out_reg_2_ ( .D(u1_fractb_s[2]), .CK(clk), .Q(fractb[2]) );
  DFF_X2 u1_fractb_out_reg_3_ ( .D(u1_fractb_s[3]), .CK(clk), .Q(fractb[3]) );
  DFF_X2 u1_fractb_out_reg_4_ ( .D(u1_fractb_s[4]), .CK(clk), .Q(fractb[4]) );
  DFF_X2 u1_fractb_out_reg_5_ ( .D(u1_fractb_s[5]), .CK(clk), .Q(fractb[5]) );
  DFF_X2 u1_fractb_out_reg_6_ ( .D(u1_fractb_s[6]), .CK(clk), .Q(fractb[6]) );
  DFF_X2 u1_fractb_out_reg_7_ ( .D(u1_fractb_s[7]), .CK(clk), .Q(fractb[7]) );
  DFF_X2 u1_fractb_out_reg_8_ ( .D(u1_fractb_s[8]), .CK(clk), .Q(fractb[8]) );
  DFF_X2 u1_fractb_out_reg_9_ ( .D(u1_fractb_s[9]), .CK(clk), .Q(fractb[9]) );
  DFF_X2 u1_fractb_out_reg_10_ ( .D(u1_fractb_s[10]), .CK(clk), .Q(fractb[10])
         );
  DFF_X2 u1_fractb_out_reg_11_ ( .D(u1_fractb_s[11]), .CK(clk), .Q(fractb[11])
         );
  DFF_X2 u1_fractb_out_reg_12_ ( .D(u1_fractb_s[12]), .CK(clk), .Q(fractb[12])
         );
  DFF_X2 u1_fractb_out_reg_13_ ( .D(u1_fractb_s[13]), .CK(clk), .Q(fractb[13])
         );
  DFF_X2 u1_fractb_out_reg_14_ ( .D(u1_fractb_s[14]), .CK(clk), .Q(fractb[14])
         );
  DFF_X2 u1_fractb_out_reg_15_ ( .D(u1_fractb_s[15]), .CK(clk), .Q(fractb[15])
         );
  DFF_X2 u1_fractb_out_reg_16_ ( .D(u1_fractb_s[16]), .CK(clk), .Q(fractb[16])
         );
  DFF_X2 u1_fractb_out_reg_17_ ( .D(u1_fractb_s[17]), .CK(clk), .Q(fractb[17])
         );
  DFF_X2 u1_fractb_out_reg_18_ ( .D(u1_fractb_s[18]), .CK(clk), .Q(fractb[18])
         );
  DFF_X2 u1_fractb_out_reg_19_ ( .D(u1_fractb_s[19]), .CK(clk), .Q(fractb[19])
         );
  DFF_X2 u1_fractb_out_reg_20_ ( .D(u1_fractb_s[20]), .CK(clk), .Q(fractb[20])
         );
  DFF_X2 u1_fractb_out_reg_21_ ( .D(u1_fractb_s[21]), .CK(clk), .Q(fractb[21])
         );
  DFF_X2 u1_fractb_out_reg_22_ ( .D(u1_fractb_s[22]), .CK(clk), .Q(fractb[22])
         );
  DFF_X2 u1_fractb_out_reg_23_ ( .D(u1_fractb_s[23]), .CK(clk), .Q(fractb[23])
         );
  DFF_X2 u1_fractb_out_reg_24_ ( .D(u1_fractb_s[24]), .CK(clk), .Q(fractb[24])
         );
  DFF_X2 u1_fractb_out_reg_25_ ( .D(u1_fractb_s[25]), .CK(clk), .Q(fractb[25])
         );
  DFF_X2 u1_fractb_out_reg_26_ ( .D(u1_fractb_s[26]), .CK(clk), .Q(fractb[26])
         );
  DFF_X2 u1_fractb_out_reg_27_ ( .D(u1_fractb_s[27]), .CK(clk), .Q(fractb[27])
         );
  DFF_X2 u1_fractb_out_reg_28_ ( .D(u1_fractb_s[28]), .CK(clk), .Q(fractb[28])
         );
  DFF_X2 u1_fractb_out_reg_29_ ( .D(u1_fractb_s[29]), .CK(clk), .Q(fractb[29])
         );
  DFF_X2 u1_fractb_out_reg_30_ ( .D(u1_fractb_s[30]), .CK(clk), .Q(fractb[30])
         );
  DFF_X2 u1_fractb_out_reg_31_ ( .D(u1_fractb_s[31]), .CK(clk), .Q(fractb[31])
         );
  DFF_X2 u1_fractb_out_reg_32_ ( .D(u1_fractb_s[32]), .CK(clk), .Q(fractb[32])
         );
  DFF_X2 u1_fractb_out_reg_33_ ( .D(u1_fractb_s[33]), .CK(clk), .Q(fractb[33])
         );
  DFF_X2 u1_fractb_out_reg_34_ ( .D(u1_fractb_s[34]), .CK(clk), .Q(fractb[34])
         );
  DFF_X2 u1_fractb_out_reg_35_ ( .D(u1_fractb_s[35]), .CK(clk), .Q(fractb[35])
         );
  DFF_X2 u1_fractb_out_reg_36_ ( .D(u1_fractb_s[36]), .CK(clk), .Q(fractb[36])
         );
  DFF_X2 u1_fractb_out_reg_37_ ( .D(u1_fractb_s[37]), .CK(clk), .Q(fractb[37])
         );
  DFF_X2 u1_fractb_out_reg_38_ ( .D(u1_fractb_s[38]), .CK(clk), .Q(fractb[38])
         );
  DFF_X2 u1_fractb_out_reg_39_ ( .D(u1_fractb_s[39]), .CK(clk), .Q(fractb[39])
         );
  DFF_X2 u1_fractb_out_reg_40_ ( .D(u1_fractb_s[40]), .CK(clk), .Q(fractb[40])
         );
  DFF_X2 u1_fractb_out_reg_41_ ( .D(u1_fractb_s[41]), .CK(clk), .Q(fractb[41])
         );
  DFF_X2 u1_fractb_out_reg_42_ ( .D(u1_fractb_s[42]), .CK(clk), .Q(fractb[42])
         );
  DFF_X2 u1_fractb_out_reg_43_ ( .D(u1_fractb_s[43]), .CK(clk), .Q(fractb[43])
         );
  DFF_X2 u1_fractb_out_reg_44_ ( .D(u1_fractb_s[44]), .CK(clk), .Q(fractb[44])
         );
  DFF_X2 u1_fractb_out_reg_45_ ( .D(u1_fractb_s[45]), .CK(clk), .Q(fractb[45])
         );
  DFF_X2 u1_fractb_out_reg_46_ ( .D(u1_fractb_s[46]), .CK(clk), .Q(fractb[46])
         );
  DFF_X2 u1_fractb_out_reg_47_ ( .D(u1_fractb_s[47]), .CK(clk), .Q(fractb[47])
         );
  DFF_X2 u1_fractb_out_reg_48_ ( .D(u1_fractb_s[48]), .CK(clk), .Q(fractb[48])
         );
  DFF_X2 u1_fractb_out_reg_49_ ( .D(u1_fractb_s[49]), .CK(clk), .Q(fractb[49])
         );
  DFF_X2 u1_fractb_out_reg_50_ ( .D(u1_fractb_s[50]), .CK(clk), .Q(fractb[50])
         );
  DFF_X2 u1_fractb_out_reg_51_ ( .D(u1_fractb_s[51]), .CK(clk), .Q(fractb[51])
         );
  DFF_X2 u1_fractb_out_reg_52_ ( .D(u1_fractb_s[52]), .CK(clk), .Q(fractb[52])
         );
  DFF_X2 u1_fractb_out_reg_53_ ( .D(u1_fractb_s[53]), .CK(clk), .Q(fractb[53])
         );
  DFF_X2 u1_fractb_out_reg_54_ ( .D(u1_fractb_s[54]), .CK(clk), .Q(fractb[54])
         );
  DFF_X2 u1_fractb_out_reg_55_ ( .D(u1_fractb_s[55]), .CK(clk), .Q(fractb[55])
         );
  DFF_X2 u1_fracta_out_reg_0_ ( .D(u1_fracta_s[0]), .CK(clk), .Q(fracta[0]) );
  DFF_X2 u1_fracta_out_reg_1_ ( .D(u1_fracta_s[1]), .CK(clk), .Q(fracta[1]) );
  DFF_X2 u1_fracta_out_reg_2_ ( .D(u1_fracta_s[2]), .CK(clk), .Q(fracta[2]) );
  DFF_X2 u1_fracta_out_reg_3_ ( .D(u1_fracta_s[3]), .CK(clk), .Q(fracta[3]) );
  DFF_X2 u1_fracta_out_reg_4_ ( .D(u1_fracta_s[4]), .CK(clk), .Q(fracta[4]) );
  DFF_X2 u1_fracta_out_reg_5_ ( .D(u1_fracta_s[5]), .CK(clk), .Q(fracta[5]) );
  DFF_X2 u1_fracta_out_reg_6_ ( .D(u1_fracta_s[6]), .CK(clk), .Q(fracta[6]) );
  DFF_X2 u1_fracta_out_reg_7_ ( .D(u1_fracta_s[7]), .CK(clk), .Q(fracta[7]) );
  DFF_X2 u1_fracta_out_reg_8_ ( .D(u1_fracta_s[8]), .CK(clk), .Q(fracta[8]) );
  DFF_X2 u1_fracta_out_reg_9_ ( .D(u1_fracta_s[9]), .CK(clk), .Q(fracta[9]) );
  DFF_X2 u1_fracta_out_reg_10_ ( .D(u1_fracta_s[10]), .CK(clk), .Q(fracta[10])
         );
  DFF_X2 u1_fracta_out_reg_11_ ( .D(u1_fracta_s[11]), .CK(clk), .Q(fracta[11])
         );
  DFF_X2 u1_fracta_out_reg_12_ ( .D(u1_fracta_s[12]), .CK(clk), .Q(fracta[12])
         );
  DFF_X2 u1_fracta_out_reg_13_ ( .D(u1_fracta_s[13]), .CK(clk), .Q(fracta[13])
         );
  DFF_X2 u1_fracta_out_reg_14_ ( .D(u1_fracta_s[14]), .CK(clk), .Q(fracta[14])
         );
  DFF_X2 u1_fracta_out_reg_15_ ( .D(u1_fracta_s[15]), .CK(clk), .Q(fracta[15])
         );
  DFF_X2 u1_fracta_out_reg_16_ ( .D(u1_fracta_s[16]), .CK(clk), .Q(fracta[16])
         );
  DFF_X2 u1_fracta_out_reg_17_ ( .D(u1_fracta_s[17]), .CK(clk), .Q(fracta[17])
         );
  DFF_X2 u1_fracta_out_reg_18_ ( .D(u1_fracta_s[18]), .CK(clk), .Q(fracta[18])
         );
  DFF_X2 u1_fracta_out_reg_19_ ( .D(u1_fracta_s[19]), .CK(clk), .Q(fracta[19])
         );
  DFF_X2 u1_fracta_out_reg_20_ ( .D(u1_fracta_s[20]), .CK(clk), .Q(fracta[20])
         );
  DFF_X2 u1_fracta_out_reg_21_ ( .D(u1_fracta_s[21]), .CK(clk), .Q(fracta[21])
         );
  DFF_X2 u1_fracta_out_reg_22_ ( .D(u1_fracta_s[22]), .CK(clk), .Q(fracta[22])
         );
  DFF_X2 u1_fracta_out_reg_23_ ( .D(u1_fracta_s[23]), .CK(clk), .Q(fracta[23])
         );
  DFF_X2 u1_fracta_out_reg_24_ ( .D(u1_fracta_s[24]), .CK(clk), .Q(fracta[24])
         );
  DFF_X2 u1_fracta_out_reg_25_ ( .D(u1_fracta_s[25]), .CK(clk), .Q(fracta[25])
         );
  DFF_X2 u1_fracta_out_reg_26_ ( .D(u1_fracta_s[26]), .CK(clk), .Q(fracta[26])
         );
  DFF_X2 u1_fracta_out_reg_27_ ( .D(u1_fracta_s[27]), .CK(clk), .Q(fracta[27])
         );
  DFF_X2 u1_fracta_out_reg_28_ ( .D(u1_fracta_s[28]), .CK(clk), .Q(fracta[28])
         );
  DFF_X2 u1_fracta_out_reg_29_ ( .D(u1_fracta_s[29]), .CK(clk), .Q(fracta[29])
         );
  DFF_X2 u1_fracta_out_reg_30_ ( .D(u1_fracta_s[30]), .CK(clk), .Q(fracta[30])
         );
  DFF_X2 u1_fracta_out_reg_31_ ( .D(u1_fracta_s[31]), .CK(clk), .Q(fracta[31])
         );
  DFF_X2 u1_fracta_out_reg_32_ ( .D(u1_fracta_s[32]), .CK(clk), .Q(fracta[32])
         );
  DFF_X2 u1_fracta_out_reg_33_ ( .D(u1_fracta_s[33]), .CK(clk), .Q(fracta[33])
         );
  DFF_X2 u1_fracta_out_reg_34_ ( .D(u1_fracta_s[34]), .CK(clk), .Q(fracta[34])
         );
  DFF_X2 u1_fracta_out_reg_35_ ( .D(u1_fracta_s[35]), .CK(clk), .Q(fracta[35])
         );
  DFF_X2 u1_fracta_out_reg_36_ ( .D(u1_fracta_s[36]), .CK(clk), .Q(fracta[36])
         );
  DFF_X2 u1_fracta_out_reg_37_ ( .D(u1_fracta_s[37]), .CK(clk), .Q(fracta[37])
         );
  DFF_X2 u1_fracta_out_reg_38_ ( .D(u1_fracta_s[38]), .CK(clk), .Q(fracta[38])
         );
  DFF_X2 u1_fracta_out_reg_39_ ( .D(u1_fracta_s[39]), .CK(clk), .Q(fracta[39])
         );
  DFF_X2 u1_fracta_out_reg_40_ ( .D(u1_fracta_s[40]), .CK(clk), .Q(fracta[40])
         );
  DFF_X2 u1_fracta_out_reg_41_ ( .D(u1_fracta_s[41]), .CK(clk), .Q(fracta[41])
         );
  DFF_X2 u1_fracta_out_reg_42_ ( .D(u1_fracta_s[42]), .CK(clk), .Q(fracta[42])
         );
  DFF_X2 u1_fracta_out_reg_43_ ( .D(u1_fracta_s[43]), .CK(clk), .Q(fracta[43])
         );
  DFF_X2 u1_fracta_out_reg_44_ ( .D(u1_fracta_s[44]), .CK(clk), .Q(fracta[44])
         );
  DFF_X2 u1_fracta_out_reg_45_ ( .D(u1_fracta_s[45]), .CK(clk), .Q(fracta[45])
         );
  DFF_X2 u1_fracta_out_reg_46_ ( .D(u1_fracta_s[46]), .CK(clk), .Q(fracta[46])
         );
  DFF_X2 u1_fracta_out_reg_47_ ( .D(u1_fracta_s[47]), .CK(clk), .Q(fracta[47])
         );
  DFF_X2 u1_fracta_out_reg_48_ ( .D(u1_fracta_s[48]), .CK(clk), .Q(fracta[48])
         );
  DFF_X2 u1_fracta_out_reg_49_ ( .D(u1_fracta_s[49]), .CK(clk), .Q(fracta[49])
         );
  DFF_X2 u1_fracta_out_reg_50_ ( .D(u1_fracta_s[50]), .CK(clk), .Q(fracta[50])
         );
  DFF_X2 u1_fracta_out_reg_51_ ( .D(u1_fracta_s[51]), .CK(clk), .Q(fracta[51])
         );
  DFF_X2 u1_fracta_out_reg_52_ ( .D(u1_fracta_s[52]), .CK(clk), .Q(fracta[52])
         );
  DFF_X2 u1_fracta_out_reg_53_ ( .D(u1_fracta_s[53]), .CK(clk), .Q(fracta[53])
         );
  DFF_X2 u1_fracta_out_reg_54_ ( .D(u1_fracta_s[54]), .CK(clk), .Q(fracta[54])
         );
  DFF_X2 u1_fracta_out_reg_55_ ( .D(u1_fracta_s[55]), .CK(clk), .Q(fracta[55])
         );
  DFF_X2 fract_out_q_reg_0_ ( .D(n6093), .CK(clk), .Q(fract_out_q[0]) );
  DFF_X2 fract_out_q_reg_1_ ( .D(n6092), .CK(clk), .Q(fract_out_q[1]) );
  DFF_X2 fract_out_q_reg_2_ ( .D(n6091), .CK(clk), .Q(fract_out_q[2]) );
  DFF_X2 fract_out_q_reg_3_ ( .D(n6090), .CK(clk), .Q(fract_out_q[3]) );
  DFF_X2 fract_out_q_reg_4_ ( .D(n6089), .CK(clk), .Q(fract_out_q[4]) );
  DFF_X2 fract_out_q_reg_5_ ( .D(n6088), .CK(clk), .Q(fract_out_q[5]) );
  DFF_X2 fract_out_q_reg_6_ ( .D(n6087), .CK(clk), .Q(fract_out_q[6]) );
  DFF_X2 fract_out_q_reg_7_ ( .D(n6086), .CK(clk), .Q(fract_out_q[7]) );
  DFF_X2 fract_out_q_reg_8_ ( .D(n6085), .CK(clk), .Q(fract_out_q[8]) );
  DFF_X2 fract_out_q_reg_9_ ( .D(n6084), .CK(clk), .Q(fract_out_q[9]) );
  DFF_X2 fract_out_q_reg_10_ ( .D(n6083), .CK(clk), .Q(fract_out_q[10]) );
  DFF_X2 fract_out_q_reg_11_ ( .D(n6082), .CK(clk), .Q(fract_out_q[11]) );
  DFF_X2 fract_out_q_reg_12_ ( .D(n6081), .CK(clk), .Q(fract_out_q[12]) );
  DFF_X2 fract_out_q_reg_13_ ( .D(n6080), .CK(clk), .Q(fract_out_q[13]) );
  DFF_X2 fract_out_q_reg_14_ ( .D(n6079), .CK(clk), .Q(fract_out_q[14]) );
  DFF_X2 fract_out_q_reg_15_ ( .D(n6078), .CK(clk), .Q(fract_out_q[15]) );
  DFF_X2 fract_out_q_reg_16_ ( .D(n6077), .CK(clk), .Q(fract_out_q[16]) );
  DFF_X2 fract_out_q_reg_17_ ( .D(n6076), .CK(clk), .Q(fract_out_q[17]) );
  DFF_X2 fract_out_q_reg_18_ ( .D(n6075), .CK(clk), .Q(fract_out_q[18]) );
  DFF_X2 fract_out_q_reg_19_ ( .D(n6074), .CK(clk), .Q(fract_out_q[19]) );
  DFF_X2 fract_out_q_reg_20_ ( .D(n6073), .CK(clk), .Q(fract_out_q[20]) );
  DFF_X2 fract_out_q_reg_21_ ( .D(n6072), .CK(clk), .Q(fract_out_q[21]) );
  DFF_X2 fract_out_q_reg_22_ ( .D(n6071), .CK(clk), .Q(fract_out_q[22]) );
  DFF_X2 fract_out_q_reg_23_ ( .D(n6070), .CK(clk), .Q(fract_out_q[23]) );
  DFF_X2 fract_out_q_reg_24_ ( .D(n6069), .CK(clk), .Q(fract_out_q[24]) );
  DFF_X2 fract_out_q_reg_25_ ( .D(n6068), .CK(clk), .Q(fract_out_q[25]) );
  DFF_X2 fract_out_q_reg_26_ ( .D(n6067), .CK(clk), .Q(fract_out_q[26]) );
  DFF_X2 fract_out_q_reg_27_ ( .D(n6066), .CK(clk), .Q(fract_out_q[27]) );
  DFF_X2 fract_out_q_reg_28_ ( .D(n6065), .CK(clk), .Q(fract_out_q[28]) );
  DFF_X2 fract_out_q_reg_29_ ( .D(n6064), .CK(clk), .Q(fract_out_q[29]) );
  DFF_X2 fract_out_q_reg_30_ ( .D(n6063), .CK(clk), .Q(fract_out_q[30]) );
  DFF_X2 fract_out_q_reg_31_ ( .D(n6062), .CK(clk), .Q(fract_out_q[31]) );
  DFF_X2 fract_out_q_reg_32_ ( .D(n6061), .CK(clk), .Q(fract_out_q[32]) );
  DFF_X2 fract_out_q_reg_33_ ( .D(n6060), .CK(clk), .Q(fract_out_q[33]) );
  DFF_X2 fract_out_q_reg_34_ ( .D(n6059), .CK(clk), .Q(fract_out_q[34]) );
  DFF_X2 fract_out_q_reg_35_ ( .D(n6058), .CK(clk), .Q(fract_out_q[35]) );
  DFF_X2 fract_out_q_reg_36_ ( .D(n6057), .CK(clk), .Q(fract_out_q[36]) );
  DFF_X2 fract_out_q_reg_37_ ( .D(n6056), .CK(clk), .Q(fract_out_q[37]) );
  DFF_X2 fract_out_q_reg_38_ ( .D(n6055), .CK(clk), .Q(fract_out_q[38]) );
  DFF_X2 fract_out_q_reg_39_ ( .D(n6054), .CK(clk), .Q(fract_out_q[39]) );
  DFF_X2 fract_out_q_reg_40_ ( .D(n6053), .CK(clk), .Q(fract_out_q[40]) );
  DFF_X2 fract_out_q_reg_41_ ( .D(n6052), .CK(clk), .Q(fract_out_q[41]) );
  DFF_X2 fract_out_q_reg_42_ ( .D(n6051), .CK(clk), .Q(fract_out_q[42]) );
  DFF_X2 fract_out_q_reg_43_ ( .D(n6050), .CK(clk), .Q(fract_out_q[43]) );
  DFF_X2 fract_out_q_reg_44_ ( .D(n6049), .CK(clk), .Q(fract_out_q[44]) );
  DFF_X2 fract_out_q_reg_45_ ( .D(n6048), .CK(clk), .Q(fract_out_q[45]) );
  DFF_X2 fract_out_q_reg_46_ ( .D(n6047), .CK(clk), .Q(fract_out_q[46]) );
  DFF_X2 fract_out_q_reg_47_ ( .D(n6046), .CK(clk), .Q(fract_out_q[47]) );
  DFF_X2 fract_out_q_reg_48_ ( .D(n6045), .CK(clk), .Q(fract_out_q[48]) );
  DFF_X2 fract_out_q_reg_49_ ( .D(n6044), .CK(clk), .Q(fract_out_q[49]) );
  DFF_X2 fract_out_q_reg_50_ ( .D(n6043), .CK(clk), .Q(fract_out_q[50]) );
  DFF_X2 fract_out_q_reg_51_ ( .D(n6042), .CK(clk), .Q(fract_out_q[51]) );
  DFF_X2 fract_out_q_reg_52_ ( .D(n6041), .CK(clk), .Q(fract_out_q[52]) );
  DFF_X2 fract_out_q_reg_53_ ( .D(n6040), .CK(clk), .Q(fract_out_q[53]) );
  DFF_X2 fract_out_q_reg_54_ ( .D(n6039), .CK(clk), .Q(fract_out_q[54]) );
  DFF_X2 fract_out_q_reg_55_ ( .D(n6038), .CK(clk), .Q(fract_out_q[55]) );
  DFF_X2 fract_out_q_reg_56_ ( .D(n6037), .CK(clk), .Q(fract_out_q[56]) );
  DFF_X2 u1_exp_dn_out_reg_0_ ( .D(u1_N52), .CK(clk), .Q(exp_fasu[0]) );
  DFF_X2 u1_exp_dn_out_reg_1_ ( .D(u1_N53), .CK(clk), .Q(exp_fasu[1]) );
  DFF_X2 u1_exp_dn_out_reg_2_ ( .D(u1_N54), .CK(clk), .Q(exp_fasu[2]) );
  DFF_X2 u1_exp_dn_out_reg_3_ ( .D(u1_N55), .CK(clk), .Q(exp_fasu[3]) );
  DFF_X2 u1_exp_dn_out_reg_4_ ( .D(u1_N56), .CK(clk), .Q(exp_fasu[4]) );
  DFF_X2 u1_exp_dn_out_reg_5_ ( .D(u1_N57), .CK(clk), .Q(exp_fasu[5]) );
  DFF_X2 u1_exp_dn_out_reg_6_ ( .D(u1_N58), .CK(clk), .Q(exp_fasu[6]) );
  DFF_X2 u1_exp_dn_out_reg_7_ ( .D(u1_N59), .CK(clk), .Q(exp_fasu[7]) );
  DFF_X2 u1_exp_dn_out_reg_8_ ( .D(u1_N60), .CK(clk), .Q(exp_fasu[8]) );
  DFF_X2 u1_exp_dn_out_reg_9_ ( .D(u1_N61), .CK(clk), .Q(exp_fasu[9]) );
  DFF_X2 u1_exp_dn_out_reg_10_ ( .D(u1_N62), .CK(clk), .Q(exp_fasu[10]) );
  DFF_X2 u2_sign_exe_reg ( .D(u2_N121), .CK(clk), .Q(sign_exe) );
  DFF_X2 sign_exe_r_reg ( .D(sign_exe), .CK(clk), .QN(n4482) );
  DFF_X2 u2_sign_reg ( .D(u2_sign_d), .CK(clk), .Q(sign_mul) );
  DFF_X2 sign_mul_r_reg ( .D(sign_mul), .CK(clk), .Q(sign_mul_r), .QN(n4491)
         );
  DFF_X2 sign_reg ( .D(N789), .CK(clk), .Q(sign), .QN(n4485) );
  DFF_X2 fract_i2f_reg_105_ ( .D(N769), .CK(clk), .Q(fract_i2f[105]) );
  DFF_X2 fract_i2f_reg_104_ ( .D(N768), .CK(clk), .Q(fract_i2f[104]) );
  DFF_X2 fract_i2f_reg_103_ ( .D(N767), .CK(clk), .Q(fract_i2f[103]) );
  DFF_X2 fract_i2f_reg_102_ ( .D(N766), .CK(clk), .Q(fract_i2f[102]) );
  DFF_X2 fract_i2f_reg_101_ ( .D(N765), .CK(clk), .Q(fract_i2f[101]) );
  DFF_X2 fract_i2f_reg_100_ ( .D(N764), .CK(clk), .Q(fract_i2f[100]) );
  DFF_X2 fract_i2f_reg_99_ ( .D(N763), .CK(clk), .Q(fract_i2f[99]) );
  DFF_X2 fract_i2f_reg_98_ ( .D(N762), .CK(clk), .Q(fract_i2f[98]) );
  DFF_X2 fract_i2f_reg_97_ ( .D(N761), .CK(clk), .Q(fract_i2f[97]) );
  DFF_X2 fract_i2f_reg_96_ ( .D(N760), .CK(clk), .Q(fract_i2f[96]) );
  DFF_X2 fract_i2f_reg_95_ ( .D(N759), .CK(clk), .Q(fract_i2f[95]) );
  DFF_X2 fract_i2f_reg_94_ ( .D(N758), .CK(clk), .Q(fract_i2f[94]) );
  DFF_X2 fract_i2f_reg_93_ ( .D(N757), .CK(clk), .Q(fract_i2f[93]) );
  DFF_X2 fract_i2f_reg_92_ ( .D(N756), .CK(clk), .Q(fract_i2f[92]) );
  DFF_X2 fract_i2f_reg_91_ ( .D(N755), .CK(clk), .Q(fract_i2f[91]) );
  DFF_X2 fract_i2f_reg_90_ ( .D(N754), .CK(clk), .Q(fract_i2f[90]) );
  DFF_X2 fract_i2f_reg_89_ ( .D(N753), .CK(clk), .Q(fract_i2f[89]) );
  DFF_X2 fract_i2f_reg_88_ ( .D(N752), .CK(clk), .Q(fract_i2f[88]) );
  DFF_X2 fract_i2f_reg_87_ ( .D(N751), .CK(clk), .Q(fract_i2f[87]) );
  DFF_X2 fract_i2f_reg_86_ ( .D(N750), .CK(clk), .Q(fract_i2f[86]) );
  DFF_X2 fract_i2f_reg_85_ ( .D(N749), .CK(clk), .Q(fract_i2f[85]) );
  DFF_X2 fract_i2f_reg_84_ ( .D(N748), .CK(clk), .Q(fract_i2f[84]) );
  DFF_X2 fract_i2f_reg_83_ ( .D(N747), .CK(clk), .Q(fract_i2f[83]) );
  DFF_X2 fract_i2f_reg_82_ ( .D(N746), .CK(clk), .Q(fract_i2f[82]) );
  DFF_X2 fract_i2f_reg_81_ ( .D(N745), .CK(clk), .Q(fract_i2f[81]) );
  DFF_X2 fract_i2f_reg_80_ ( .D(N744), .CK(clk), .Q(fract_i2f[80]) );
  DFF_X2 fract_i2f_reg_79_ ( .D(N743), .CK(clk), .Q(fract_i2f[79]) );
  DFF_X2 fract_i2f_reg_78_ ( .D(N742), .CK(clk), .Q(fract_i2f[78]) );
  DFF_X2 fract_i2f_reg_77_ ( .D(N741), .CK(clk), .Q(fract_i2f[77]) );
  DFF_X2 fract_i2f_reg_76_ ( .D(N740), .CK(clk), .Q(fract_i2f[76]) );
  DFF_X2 fract_i2f_reg_75_ ( .D(N739), .CK(clk), .Q(fract_i2f[75]) );
  DFF_X2 fract_i2f_reg_74_ ( .D(N738), .CK(clk), .Q(fract_i2f[74]) );
  DFF_X2 fract_i2f_reg_73_ ( .D(N737), .CK(clk), .Q(fract_i2f[73]) );
  DFF_X2 fract_i2f_reg_72_ ( .D(N736), .CK(clk), .Q(fract_i2f[72]) );
  DFF_X2 fract_i2f_reg_71_ ( .D(N735), .CK(clk), .Q(fract_i2f[71]) );
  DFF_X2 fract_i2f_reg_70_ ( .D(N734), .CK(clk), .Q(fract_i2f[70]) );
  DFF_X2 fract_i2f_reg_69_ ( .D(N733), .CK(clk), .Q(fract_i2f[69]) );
  DFF_X2 fract_i2f_reg_68_ ( .D(N732), .CK(clk), .Q(fract_i2f[68]) );
  DFF_X2 fract_i2f_reg_67_ ( .D(N731), .CK(clk), .Q(fract_i2f[67]) );
  DFF_X2 fract_i2f_reg_66_ ( .D(N730), .CK(clk), .Q(fract_i2f[66]) );
  DFF_X2 fract_i2f_reg_65_ ( .D(N729), .CK(clk), .Q(fract_i2f[65]) );
  DFF_X2 fract_i2f_reg_64_ ( .D(N728), .CK(clk), .Q(fract_i2f[64]) );
  DFF_X2 fract_i2f_reg_63_ ( .D(N727), .CK(clk), .Q(fract_i2f[63]) );
  DFF_X2 fract_i2f_reg_62_ ( .D(N726), .CK(clk), .Q(fract_i2f[62]) );
  DFF_X2 fract_i2f_reg_61_ ( .D(N725), .CK(clk), .Q(fract_i2f[61]) );
  DFF_X2 fract_i2f_reg_60_ ( .D(N724), .CK(clk), .Q(fract_i2f[60]) );
  DFF_X2 fract_i2f_reg_59_ ( .D(N723), .CK(clk), .Q(fract_i2f[59]) );
  DFF_X2 fract_i2f_reg_58_ ( .D(N722), .CK(clk), .Q(fract_i2f[58]) );
  DFF_X2 fract_i2f_reg_57_ ( .D(N721), .CK(clk), .Q(fract_i2f[57]) );
  DFF_X2 fract_i2f_reg_56_ ( .D(N720), .CK(clk), .Q(fract_i2f[56]) );
  DFF_X2 fract_i2f_reg_55_ ( .D(N719), .CK(clk), .Q(fract_i2f[55]) );
  DFF_X2 fract_i2f_reg_54_ ( .D(N718), .CK(clk), .Q(fract_i2f[54]) );
  DFF_X2 fract_i2f_reg_53_ ( .D(N717), .CK(clk), .Q(fract_i2f[53]) );
  DFF_X2 fract_i2f_reg_52_ ( .D(N716), .CK(clk), .Q(fract_i2f[52]) );
  DFF_X2 fract_i2f_reg_51_ ( .D(N715), .CK(clk), .Q(fract_i2f[51]) );
  DFF_X2 fract_i2f_reg_50_ ( .D(N714), .CK(clk), .Q(fract_i2f[50]) );
  DFF_X2 fract_i2f_reg_49_ ( .D(N713), .CK(clk), .Q(fract_i2f[49]) );
  DFF_X2 fract_i2f_reg_48_ ( .D(N712), .CK(clk), .Q(fract_i2f[48]) );
  DFF_X2 fract_i2f_reg_47_ ( .D(N711), .CK(clk), .Q(fract_i2f[47]) );
  DFF_X2 fract_i2f_reg_46_ ( .D(N710), .CK(clk), .Q(fract_i2f[46]) );
  DFF_X2 fract_i2f_reg_45_ ( .D(n5913), .CK(clk), .Q(fract_i2f[45]) );
  DFF_X2 fract_i2f_reg_44_ ( .D(n5914), .CK(clk), .Q(fract_i2f[44]) );
  DFF_X2 fract_i2f_reg_43_ ( .D(n5915), .CK(clk), .Q(fract_i2f[43]) );
  DFF_X2 fract_i2f_reg_42_ ( .D(n5916), .CK(clk), .Q(fract_i2f[42]) );
  DFF_X2 fract_i2f_reg_41_ ( .D(n5917), .CK(clk), .Q(fract_i2f[41]) );
  DFF_X2 fract_i2f_reg_40_ ( .D(n5918), .CK(clk), .Q(fract_i2f[40]) );
  DFF_X2 fract_i2f_reg_39_ ( .D(n5919), .CK(clk), .Q(fract_i2f[39]) );
  DFF_X2 fract_i2f_reg_38_ ( .D(n5920), .CK(clk), .Q(fract_i2f[38]) );
  DFF_X2 fract_i2f_reg_37_ ( .D(n5921), .CK(clk), .Q(fract_i2f[37]) );
  DFF_X2 fract_i2f_reg_36_ ( .D(n5922), .CK(clk), .Q(fract_i2f[36]) );
  DFF_X2 fract_i2f_reg_35_ ( .D(n5923), .CK(clk), .Q(fract_i2f[35]) );
  DFF_X2 fract_i2f_reg_34_ ( .D(n5924), .CK(clk), .Q(fract_i2f[34]) );
  DFF_X2 fract_i2f_reg_33_ ( .D(n5925), .CK(clk), .Q(fract_i2f[33]) );
  DFF_X2 fract_i2f_reg_32_ ( .D(n5926), .CK(clk), .Q(fract_i2f[32]) );
  DFF_X2 fract_i2f_reg_31_ ( .D(n5927), .CK(clk), .Q(fract_i2f[31]) );
  DFF_X2 fract_i2f_reg_30_ ( .D(n5928), .CK(clk), .Q(fract_i2f[30]) );
  DFF_X2 fract_i2f_reg_29_ ( .D(n5929), .CK(clk), .Q(fract_i2f[29]) );
  DFF_X2 fract_i2f_reg_28_ ( .D(n5930), .CK(clk), .Q(fract_i2f[28]) );
  DFF_X2 fract_i2f_reg_27_ ( .D(n5931), .CK(clk), .Q(fract_i2f[27]) );
  DFF_X2 fract_i2f_reg_26_ ( .D(n5932), .CK(clk), .Q(fract_i2f[26]) );
  DFF_X2 fract_i2f_reg_25_ ( .D(n5933), .CK(clk), .Q(fract_i2f[25]) );
  DFF_X2 fract_i2f_reg_24_ ( .D(n5934), .CK(clk), .Q(fract_i2f[24]) );
  DFF_X2 fract_i2f_reg_23_ ( .D(n5935), .CK(clk), .Q(fract_i2f[23]) );
  DFF_X2 fract_i2f_reg_22_ ( .D(n5936), .CK(clk), .Q(fract_i2f[22]) );
  DFF_X2 fract_i2f_reg_21_ ( .D(n5937), .CK(clk), .Q(fract_i2f[21]) );
  DFF_X2 fract_i2f_reg_20_ ( .D(n5938), .CK(clk), .Q(fract_i2f[20]) );
  DFF_X2 fract_i2f_reg_19_ ( .D(n5939), .CK(clk), .Q(fract_i2f[19]) );
  DFF_X2 fract_i2f_reg_18_ ( .D(n5940), .CK(clk), .Q(fract_i2f[18]) );
  DFF_X2 fract_i2f_reg_17_ ( .D(n5941), .CK(clk), .Q(fract_i2f[17]) );
  DFF_X2 fract_i2f_reg_16_ ( .D(n5942), .CK(clk), .Q(fract_i2f[16]) );
  DFF_X2 fract_i2f_reg_15_ ( .D(n5943), .CK(clk), .Q(fract_i2f[15]) );
  DFF_X2 fract_i2f_reg_14_ ( .D(n5944), .CK(clk), .Q(fract_i2f[14]) );
  DFF_X2 fract_i2f_reg_13_ ( .D(n5945), .CK(clk), .Q(fract_i2f[13]) );
  DFF_X2 fract_i2f_reg_12_ ( .D(n5946), .CK(clk), .Q(fract_i2f[12]) );
  DFF_X2 fract_i2f_reg_11_ ( .D(n5947), .CK(clk), .Q(fract_i2f[11]) );
  DFF_X2 fract_i2f_reg_10_ ( .D(n5948), .CK(clk), .Q(fract_i2f[10]) );
  DFF_X2 fract_i2f_reg_9_ ( .D(n5949), .CK(clk), .Q(fract_i2f[9]) );
  DFF_X2 fract_i2f_reg_8_ ( .D(n5950), .CK(clk), .Q(fract_i2f[8]) );
  DFF_X2 fract_i2f_reg_7_ ( .D(n5951), .CK(clk), .Q(fract_i2f[7]) );
  DFF_X2 fract_i2f_reg_6_ ( .D(n5952), .CK(clk), .Q(fract_i2f[6]) );
  DFF_X2 fract_i2f_reg_5_ ( .D(n5953), .CK(clk), .Q(fract_i2f[5]) );
  DFF_X2 fract_i2f_reg_4_ ( .D(n5954), .CK(clk), .Q(fract_i2f[4]) );
  DFF_X2 fract_i2f_reg_3_ ( .D(n5955), .CK(clk), .Q(fract_i2f[3]) );
  DFF_X2 fract_i2f_reg_2_ ( .D(n5956), .CK(clk), .Q(fract_i2f[2]) );
  DFF_X2 fract_i2f_reg_1_ ( .D(n5957), .CK(clk), .Q(fract_i2f[1]) );
  DFF_X2 fract_i2f_reg_0_ ( .D(n6311), .CK(clk), .Q(fract_i2f[0]) );
  DFF_X2 u2_inf_reg ( .D(u2_N114), .CK(clk), .Q(inf_mul) );
  DFF_X2 inf_mul_r_reg ( .D(inf_mul), .CK(clk), .Q(inf_mul_r) );
  DFF_X2 u2_underflow_reg_0_ ( .D(u2_underflow_d[0]), .CK(clk), .Q(
        underflow_fmul_d[0]) );
  DFF_X2 underflow_fmul_r_reg_0_ ( .D(underflow_fmul_d[0]), .CK(clk), .Q(
        underflow_fmul_r[0]) );
  DFF_X2 u2_underflow_reg_1_ ( .D(u2_underflow_d[1]), .CK(clk), .Q(
        underflow_fmul_d[1]) );
  DFF_X2 underflow_fmul_r_reg_1_ ( .D(underflow_fmul_d[1]), .CK(clk), .Q(
        underflow_fmul_r[1]) );
  DFF_X2 u2_underflow_reg_2_ ( .D(u2_underflow_d[2]), .CK(clk), .Q(
        underflow_fmul_d[2]) );
  DFF_X2 underflow_fmul_r_reg_2_ ( .D(underflow_fmul_d[2]), .CK(clk), .Q(
        underflow_fmul_r[2]) );
  DFF_X2 u2_exp_ovf_reg_0_ ( .D(u2_exp_ovf_d_0_), .CK(clk), .Q(exp_ovf[0]) );
  DFF_X2 exp_ovf_r_reg_0_ ( .D(exp_ovf[0]), .CK(clk), .Q(exp_ovf_r[0]), .QN(
        n4356) );
  DFF_X2 u2_exp_ovf_reg_1_ ( .D(u2_exp_ovf_d_1_), .CK(clk), .Q(exp_ovf[1]) );
  DFF_X2 exp_ovf_r_reg_1_ ( .D(exp_ovf[1]), .CK(clk), .Q(exp_ovf_r[1]), .QN(
        n4452) );
  DFF_X2 u2_exp_out_reg_0_ ( .D(u2_N76), .CK(clk), .QN(n4383) );
  DFF_X2 exp_r_reg_0_ ( .D(N327), .CK(clk), .QN(n4349) );
  DFF_X2 u2_exp_out_reg_1_ ( .D(u2_N77), .CK(clk), .QN(n4487) );
  DFF_X2 exp_r_reg_1_ ( .D(N328), .CK(clk), .Q(exp_r[1]), .QN(n4314) );
  DFF_X2 u2_exp_out_reg_2_ ( .D(u2_N78), .CK(clk), .Q(exp_mul[2]), .QN(n4539)
         );
  DFF_X2 exp_r_reg_2_ ( .D(N329), .CK(clk), .Q(n4315), .QN(n4438) );
  DFF_X2 u2_exp_out_reg_3_ ( .D(u2_N79), .CK(clk), .Q(exp_mul[3]), .QN(n4538)
         );
  DFF_X2 exp_r_reg_3_ ( .D(N330), .CK(clk), .Q(exp_r[3]), .QN(n4316) );
  DFF_X2 u2_exp_out_reg_4_ ( .D(u2_N80), .CK(clk), .Q(exp_mul[4]), .QN(n4537)
         );
  DFF_X2 exp_r_reg_4_ ( .D(N331), .CK(clk), .Q(n4282), .QN(n4299) );
  DFF_X2 u2_exp_out_reg_5_ ( .D(u2_N81), .CK(clk), .Q(exp_mul[5]), .QN(n4535)
         );
  DFF_X2 exp_r_reg_5_ ( .D(N332), .CK(clk), .Q(n4290), .QN(n4347) );
  DFF_X2 u2_exp_out_reg_6_ ( .D(u2_N82), .CK(clk), .Q(exp_mul[6]), .QN(n4536)
         );
  DFF_X2 exp_r_reg_6_ ( .D(N333), .CK(clk), .Q(exp_r[6]), .QN(n4317) );
  DFF_X2 u2_exp_out_reg_7_ ( .D(u2_N83), .CK(clk), .Q(exp_mul[7]), .QN(n4534)
         );
  DFF_X2 exp_r_reg_7_ ( .D(N334), .CK(clk), .Q(n4281), .QN(n4348) );
  DFF_X2 u2_exp_out_reg_8_ ( .D(u2_N84), .CK(clk), .QN(n4489) );
  DFF_X2 exp_r_reg_8_ ( .D(N335), .CK(clk), .Q(n4353), .QN(n4439) );
  DFF_X2 u2_exp_out_reg_9_ ( .D(u2_N85), .CK(clk), .QN(n4384) );
  DFF_X2 exp_r_reg_9_ ( .D(N336), .CK(clk), .Q(n4289), .QN(n4350) );
  DFF_X2 u2_exp_out_reg_10_ ( .D(u2_N86), .CK(clk), .QN(n4330) );
  DFF_X2 inf_mul2_reg ( .D(N923), .CK(clk), .Q(inf_mul2) );
  DFF_X2 exp_r_reg_10_ ( .D(N337), .CK(clk), .Q(n4352), .QN(n4440) );
  DFF_X2 u5_prod1_reg_0_ ( .D(u5_N0), .CK(clk), .Q(u5_prod1[0]) );
  DFF_X2 u5_prod_reg_0_ ( .D(u5_prod1[0]), .CK(clk), .Q(prod[0]) );
  DFF_X2 u5_prod1_reg_1_ ( .D(u5_N1), .CK(clk), .Q(u5_prod1[1]) );
  DFF_X2 u5_prod_reg_1_ ( .D(u5_prod1[1]), .CK(clk), .Q(prod[1]) );
  DFF_X2 u5_prod1_reg_2_ ( .D(u5_N2), .CK(clk), .Q(u5_prod1[2]) );
  DFF_X2 u5_prod_reg_2_ ( .D(u5_prod1[2]), .CK(clk), .Q(prod[2]) );
  DFF_X2 u5_prod1_reg_3_ ( .D(u5_N3), .CK(clk), .Q(u5_prod1[3]) );
  DFF_X2 u5_prod_reg_3_ ( .D(u5_prod1[3]), .CK(clk), .Q(prod[3]) );
  DFF_X2 u5_prod1_reg_4_ ( .D(u5_N4), .CK(clk), .Q(u5_prod1[4]) );
  DFF_X2 u5_prod_reg_4_ ( .D(u5_prod1[4]), .CK(clk), .Q(prod[4]) );
  DFF_X2 u5_prod1_reg_5_ ( .D(u5_N5), .CK(clk), .Q(u5_prod1[5]) );
  DFF_X2 u5_prod_reg_5_ ( .D(u5_prod1[5]), .CK(clk), .Q(prod[5]) );
  DFF_X2 u5_prod1_reg_6_ ( .D(u5_N6), .CK(clk), .Q(u5_prod1[6]) );
  DFF_X2 u5_prod_reg_6_ ( .D(u5_prod1[6]), .CK(clk), .Q(prod[6]) );
  DFF_X2 u5_prod1_reg_7_ ( .D(u5_N7), .CK(clk), .Q(u5_prod1[7]) );
  DFF_X2 u5_prod_reg_7_ ( .D(u5_prod1[7]), .CK(clk), .Q(prod[7]) );
  DFF_X2 u5_prod1_reg_8_ ( .D(u5_N8), .CK(clk), .Q(u5_prod1[8]) );
  DFF_X2 u5_prod_reg_8_ ( .D(u5_prod1[8]), .CK(clk), .Q(prod[8]) );
  DFF_X2 u5_prod1_reg_9_ ( .D(u5_N9), .CK(clk), .Q(u5_prod1[9]) );
  DFF_X2 u5_prod_reg_9_ ( .D(u5_prod1[9]), .CK(clk), .Q(prod[9]) );
  DFF_X2 u5_prod1_reg_10_ ( .D(u5_N10), .CK(clk), .Q(u5_prod1[10]) );
  DFF_X2 u5_prod_reg_10_ ( .D(u5_prod1[10]), .CK(clk), .Q(prod[10]) );
  DFF_X2 u5_prod1_reg_11_ ( .D(u5_N11), .CK(clk), .Q(u5_prod1[11]) );
  DFF_X2 u5_prod_reg_11_ ( .D(u5_prod1[11]), .CK(clk), .Q(prod[11]) );
  DFF_X2 u5_prod1_reg_12_ ( .D(u5_N12), .CK(clk), .Q(u5_prod1[12]) );
  DFF_X2 u5_prod_reg_12_ ( .D(u5_prod1[12]), .CK(clk), .Q(prod[12]) );
  DFF_X2 u5_prod1_reg_13_ ( .D(u5_N13), .CK(clk), .Q(u5_prod1[13]) );
  DFF_X2 u5_prod_reg_13_ ( .D(u5_prod1[13]), .CK(clk), .Q(prod[13]) );
  DFF_X2 u5_prod1_reg_14_ ( .D(u5_N14), .CK(clk), .Q(u5_prod1[14]) );
  DFF_X2 u5_prod_reg_14_ ( .D(u5_prod1[14]), .CK(clk), .Q(prod[14]) );
  DFF_X2 u5_prod1_reg_15_ ( .D(u5_N15), .CK(clk), .Q(u5_prod1[15]) );
  DFF_X2 u5_prod_reg_15_ ( .D(u5_prod1[15]), .CK(clk), .Q(prod[15]) );
  DFF_X2 u5_prod1_reg_16_ ( .D(u5_N16), .CK(clk), .Q(u5_prod1[16]) );
  DFF_X2 u5_prod_reg_16_ ( .D(u5_prod1[16]), .CK(clk), .Q(prod[16]) );
  DFF_X2 u5_prod1_reg_17_ ( .D(u5_N17), .CK(clk), .Q(u5_prod1[17]) );
  DFF_X2 u5_prod_reg_17_ ( .D(u5_prod1[17]), .CK(clk), .Q(prod[17]) );
  DFF_X2 u5_prod1_reg_18_ ( .D(u5_N18), .CK(clk), .Q(u5_prod1[18]) );
  DFF_X2 u5_prod_reg_18_ ( .D(u5_prod1[18]), .CK(clk), .Q(prod[18]) );
  DFF_X2 u5_prod1_reg_19_ ( .D(u5_N19), .CK(clk), .Q(u5_prod1[19]) );
  DFF_X2 u5_prod_reg_19_ ( .D(u5_prod1[19]), .CK(clk), .Q(prod[19]) );
  DFF_X2 u5_prod1_reg_20_ ( .D(u5_N20), .CK(clk), .Q(u5_prod1[20]) );
  DFF_X2 u5_prod_reg_20_ ( .D(u5_prod1[20]), .CK(clk), .Q(prod[20]) );
  DFF_X2 u5_prod1_reg_21_ ( .D(u5_N21), .CK(clk), .Q(u5_prod1[21]) );
  DFF_X2 u5_prod_reg_21_ ( .D(u5_prod1[21]), .CK(clk), .Q(prod[21]) );
  DFF_X2 u5_prod1_reg_22_ ( .D(u5_N22), .CK(clk), .Q(u5_prod1[22]) );
  DFF_X2 u5_prod_reg_22_ ( .D(u5_prod1[22]), .CK(clk), .Q(prod[22]) );
  DFF_X2 u5_prod1_reg_23_ ( .D(u5_N23), .CK(clk), .Q(u5_prod1[23]) );
  DFF_X2 u5_prod_reg_23_ ( .D(u5_prod1[23]), .CK(clk), .Q(prod[23]) );
  DFF_X2 u5_prod1_reg_24_ ( .D(u5_N24), .CK(clk), .Q(u5_prod1[24]) );
  DFF_X2 u5_prod_reg_24_ ( .D(u5_prod1[24]), .CK(clk), .Q(prod[24]) );
  DFF_X2 u5_prod1_reg_25_ ( .D(u5_N25), .CK(clk), .Q(u5_prod1[25]) );
  DFF_X2 u5_prod_reg_25_ ( .D(u5_prod1[25]), .CK(clk), .Q(prod[25]) );
  DFF_X2 u5_prod1_reg_26_ ( .D(u5_N26), .CK(clk), .Q(u5_prod1[26]) );
  DFF_X2 u5_prod_reg_26_ ( .D(u5_prod1[26]), .CK(clk), .Q(prod[26]) );
  DFF_X2 u5_prod1_reg_27_ ( .D(u5_N27), .CK(clk), .Q(u5_prod1[27]) );
  DFF_X2 u5_prod_reg_27_ ( .D(u5_prod1[27]), .CK(clk), .Q(prod[27]) );
  DFF_X2 u5_prod1_reg_28_ ( .D(u5_N28), .CK(clk), .Q(u5_prod1[28]) );
  DFF_X2 u5_prod_reg_28_ ( .D(u5_prod1[28]), .CK(clk), .Q(prod[28]) );
  DFF_X2 u5_prod1_reg_29_ ( .D(u5_N29), .CK(clk), .Q(u5_prod1[29]) );
  DFF_X2 u5_prod_reg_29_ ( .D(u5_prod1[29]), .CK(clk), .Q(prod[29]) );
  DFF_X2 u5_prod1_reg_30_ ( .D(u5_N30), .CK(clk), .Q(u5_prod1[30]) );
  DFF_X2 u5_prod_reg_30_ ( .D(u5_prod1[30]), .CK(clk), .Q(prod[30]) );
  DFF_X2 u5_prod1_reg_31_ ( .D(u5_N31), .CK(clk), .Q(u5_prod1[31]) );
  DFF_X2 u5_prod_reg_31_ ( .D(u5_prod1[31]), .CK(clk), .Q(prod[31]) );
  DFF_X2 u5_prod1_reg_32_ ( .D(u5_N32), .CK(clk), .Q(u5_prod1[32]) );
  DFF_X2 u5_prod_reg_32_ ( .D(u5_prod1[32]), .CK(clk), .Q(prod[32]) );
  DFF_X2 u5_prod1_reg_33_ ( .D(u5_N33), .CK(clk), .Q(u5_prod1[33]) );
  DFF_X2 u5_prod_reg_33_ ( .D(u5_prod1[33]), .CK(clk), .Q(prod[33]) );
  DFF_X2 u5_prod1_reg_34_ ( .D(u5_N34), .CK(clk), .Q(u5_prod1[34]) );
  DFF_X2 u5_prod_reg_34_ ( .D(u5_prod1[34]), .CK(clk), .Q(prod[34]) );
  DFF_X2 u5_prod1_reg_35_ ( .D(u5_N35), .CK(clk), .Q(u5_prod1[35]) );
  DFF_X2 u5_prod_reg_35_ ( .D(u5_prod1[35]), .CK(clk), .Q(prod[35]) );
  DFF_X2 u5_prod1_reg_36_ ( .D(u5_N36), .CK(clk), .Q(u5_prod1[36]) );
  DFF_X2 u5_prod_reg_36_ ( .D(u5_prod1[36]), .CK(clk), .Q(prod[36]) );
  DFF_X2 u5_prod1_reg_37_ ( .D(u5_N37), .CK(clk), .Q(u5_prod1[37]) );
  DFF_X2 u5_prod_reg_37_ ( .D(u5_prod1[37]), .CK(clk), .Q(prod[37]) );
  DFF_X2 u5_prod1_reg_38_ ( .D(u5_N38), .CK(clk), .Q(u5_prod1[38]) );
  DFF_X2 u5_prod_reg_38_ ( .D(u5_prod1[38]), .CK(clk), .Q(prod[38]) );
  DFF_X2 u5_prod1_reg_39_ ( .D(u5_N39), .CK(clk), .Q(u5_prod1[39]) );
  DFF_X2 u5_prod_reg_39_ ( .D(u5_prod1[39]), .CK(clk), .Q(prod[39]) );
  DFF_X2 u5_prod1_reg_40_ ( .D(u5_N40), .CK(clk), .Q(u5_prod1[40]) );
  DFF_X2 u5_prod_reg_40_ ( .D(u5_prod1[40]), .CK(clk), .Q(prod[40]) );
  DFF_X2 u5_prod1_reg_41_ ( .D(u5_N41), .CK(clk), .Q(u5_prod1[41]) );
  DFF_X2 u5_prod_reg_41_ ( .D(u5_prod1[41]), .CK(clk), .Q(prod[41]) );
  DFF_X2 u5_prod1_reg_42_ ( .D(u5_N42), .CK(clk), .Q(u5_prod1[42]) );
  DFF_X2 u5_prod_reg_42_ ( .D(u5_prod1[42]), .CK(clk), .Q(prod[42]) );
  DFF_X2 u5_prod1_reg_43_ ( .D(u5_N43), .CK(clk), .Q(u5_prod1[43]) );
  DFF_X2 u5_prod_reg_43_ ( .D(u5_prod1[43]), .CK(clk), .Q(prod[43]) );
  DFF_X2 u5_prod1_reg_44_ ( .D(u5_N44), .CK(clk), .Q(u5_prod1[44]) );
  DFF_X2 u5_prod_reg_44_ ( .D(u5_prod1[44]), .CK(clk), .Q(prod[44]) );
  DFF_X2 u5_prod1_reg_45_ ( .D(u5_N45), .CK(clk), .Q(u5_prod1[45]) );
  DFF_X2 u5_prod_reg_45_ ( .D(u5_prod1[45]), .CK(clk), .Q(prod[45]) );
  DFF_X2 u5_prod1_reg_46_ ( .D(u5_N46), .CK(clk), .Q(u5_prod1[46]) );
  DFF_X2 u5_prod_reg_46_ ( .D(u5_prod1[46]), .CK(clk), .Q(prod[46]) );
  DFF_X2 u5_prod1_reg_47_ ( .D(u5_N47), .CK(clk), .Q(u5_prod1[47]) );
  DFF_X2 u5_prod_reg_47_ ( .D(u5_prod1[47]), .CK(clk), .Q(prod[47]) );
  DFF_X2 u5_prod1_reg_48_ ( .D(u5_N48), .CK(clk), .Q(u5_prod1[48]) );
  DFF_X2 u5_prod_reg_48_ ( .D(u5_prod1[48]), .CK(clk), .Q(prod[48]) );
  DFF_X2 u5_prod1_reg_49_ ( .D(u5_N49), .CK(clk), .Q(u5_prod1[49]) );
  DFF_X2 u5_prod_reg_49_ ( .D(u5_prod1[49]), .CK(clk), .Q(prod[49]) );
  DFF_X2 u5_prod1_reg_50_ ( .D(u5_N50), .CK(clk), .Q(u5_prod1[50]) );
  DFF_X2 u5_prod_reg_50_ ( .D(u5_prod1[50]), .CK(clk), .Q(prod[50]), .QN(n4434) );
  DFF_X2 u5_prod1_reg_51_ ( .D(u5_N51), .CK(clk), .Q(u5_prod1[51]) );
  DFF_X2 u5_prod_reg_51_ ( .D(u5_prod1[51]), .CK(clk), .Q(prod[51]), .QN(n4432) );
  DFF_X2 u5_prod1_reg_52_ ( .D(u5_N52), .CK(clk), .Q(u5_prod1[52]) );
  DFF_X2 u5_prod_reg_52_ ( .D(u5_prod1[52]), .CK(clk), .Q(prod[52]), .QN(n4429) );
  DFF_X2 u5_prod1_reg_53_ ( .D(u5_N53), .CK(clk), .Q(u5_prod1[53]) );
  DFF_X2 u5_prod_reg_53_ ( .D(u5_prod1[53]), .CK(clk), .Q(prod[53]), .QN(n4410) );
  DFF_X2 u5_prod1_reg_54_ ( .D(u5_N54), .CK(clk), .Q(u5_prod1[54]) );
  DFF_X2 u5_prod_reg_54_ ( .D(u5_prod1[54]), .CK(clk), .Q(prod[54]), .QN(n4419) );
  DFF_X2 u5_prod1_reg_55_ ( .D(u5_N55), .CK(clk), .Q(u5_prod1[55]) );
  DFF_X2 u5_prod_reg_55_ ( .D(u5_prod1[55]), .CK(clk), .QN(n4310) );
  DFF_X2 u5_prod1_reg_56_ ( .D(u5_N56), .CK(clk), .Q(u5_prod1[56]) );
  DFF_X2 u5_prod_reg_56_ ( .D(u5_prod1[56]), .CK(clk), .QN(n4401) );
  DFF_X2 u5_prod1_reg_57_ ( .D(u5_N57), .CK(clk), .Q(u5_prod1[57]) );
  DFF_X2 u5_prod_reg_57_ ( .D(u5_prod1[57]), .CK(clk), .QN(n4341) );
  DFF_X2 u5_prod1_reg_58_ ( .D(u5_N58), .CK(clk), .Q(u5_prod1[58]) );
  DFF_X2 u5_prod_reg_58_ ( .D(u5_prod1[58]), .CK(clk), .Q(prod[58]), .QN(n4430) );
  DFF_X2 u5_prod1_reg_59_ ( .D(u5_N59), .CK(clk), .Q(u5_prod1[59]) );
  DFF_X2 u5_prod_reg_59_ ( .D(u5_prod1[59]), .CK(clk), .Q(prod[59]), .QN(n4413) );
  DFF_X2 u5_prod1_reg_60_ ( .D(u5_N60), .CK(clk), .Q(u5_prod1[60]) );
  DFF_X2 u5_prod_reg_60_ ( .D(u5_prod1[60]), .CK(clk), .QN(n4346) );
  DFF_X2 u5_prod1_reg_61_ ( .D(u5_N61), .CK(clk), .Q(u5_prod1[61]) );
  DFF_X2 u5_prod_reg_61_ ( .D(u5_prod1[61]), .CK(clk), .QN(n4406) );
  DFF_X2 u5_prod1_reg_62_ ( .D(u5_N62), .CK(clk), .Q(u5_prod1[62]) );
  DFF_X2 u5_prod_reg_62_ ( .D(u5_prod1[62]), .CK(clk), .QN(n4312) );
  DFF_X2 u5_prod1_reg_63_ ( .D(u5_N63), .CK(clk), .Q(u5_prod1[63]) );
  DFF_X2 u5_prod_reg_63_ ( .D(u5_prod1[63]), .CK(clk), .QN(n4297) );
  DFF_X2 u5_prod1_reg_64_ ( .D(u5_N64), .CK(clk), .Q(u5_prod1[64]) );
  DFF_X2 u5_prod_reg_64_ ( .D(u5_prod1[64]), .CK(clk), .Q(prod[64]), .QN(n4428) );
  DFF_X2 u5_prod1_reg_65_ ( .D(u5_N65), .CK(clk), .Q(u5_prod1[65]) );
  DFF_X2 u5_prod_reg_65_ ( .D(u5_prod1[65]), .CK(clk), .Q(prod[65]), .QN(n4414) );
  DFF_X2 u5_prod1_reg_66_ ( .D(u5_N66), .CK(clk), .Q(u5_prod1[66]) );
  DFF_X2 u5_prod_reg_66_ ( .D(u5_prod1[66]), .CK(clk), .Q(prod[66]), .QN(n4423) );
  DFF_X2 u5_prod1_reg_67_ ( .D(u5_N67), .CK(clk), .Q(u5_prod1[67]) );
  DFF_X2 u5_prod_reg_67_ ( .D(u5_prod1[67]), .CK(clk), .QN(n4311) );
  DFF_X2 u5_prod1_reg_68_ ( .D(u5_N68), .CK(clk), .Q(u5_prod1[68]) );
  DFF_X2 u5_prod_reg_68_ ( .D(u5_prod1[68]), .CK(clk), .QN(n4402) );
  DFF_X2 u5_prod1_reg_69_ ( .D(u5_N69), .CK(clk), .Q(u5_prod1[69]) );
  DFF_X2 u5_prod_reg_69_ ( .D(u5_prod1[69]), .CK(clk), .QN(n4342) );
  DFF_X2 u5_prod1_reg_70_ ( .D(u5_N70), .CK(clk), .Q(u5_prod1[70]) );
  DFF_X2 u5_prod_reg_70_ ( .D(u5_prod1[70]), .CK(clk), .Q(prod[70]), .QN(n4415) );
  DFF_X2 u5_prod1_reg_71_ ( .D(u5_N71), .CK(clk), .Q(u5_prod1[71]) );
  DFF_X2 u5_prod_reg_71_ ( .D(u5_prod1[71]), .CK(clk), .Q(prod[71]), .QN(n4422) );
  DFF_X2 u5_prod1_reg_72_ ( .D(u5_N72), .CK(clk), .Q(u5_prod1[72]) );
  DFF_X2 u5_prod_reg_72_ ( .D(u5_prod1[72]), .CK(clk), .QN(n4313) );
  DFF_X2 u5_prod1_reg_73_ ( .D(u5_N73), .CK(clk), .Q(u5_prod1[73]) );
  DFF_X2 u5_prod_reg_73_ ( .D(u5_prod1[73]), .CK(clk), .QN(n4407) );
  DFF_X2 u5_prod1_reg_74_ ( .D(u5_N74), .CK(clk), .Q(u5_prod1[74]) );
  DFF_X2 u5_prod_reg_74_ ( .D(u5_prod1[74]), .CK(clk), .QN(n4298) );
  DFF_X2 u5_prod1_reg_75_ ( .D(u5_N75), .CK(clk), .Q(u5_prod1[75]) );
  DFF_X2 u5_prod_reg_75_ ( .D(u5_prod1[75]), .CK(clk), .QN(n4343) );
  DFF_X2 u5_prod1_reg_76_ ( .D(u5_N76), .CK(clk), .Q(u5_prod1[76]) );
  DFF_X2 u5_prod_reg_76_ ( .D(u5_prod1[76]), .CK(clk), .Q(prod[76]), .QN(n4426) );
  DFF_X2 u5_prod1_reg_77_ ( .D(u5_N77), .CK(clk), .Q(u5_prod1[77]) );
  DFF_X2 u5_prod_reg_77_ ( .D(u5_prod1[77]), .CK(clk), .Q(prod[77]), .QN(n4412) );
  DFF_X2 u5_prod1_reg_78_ ( .D(u5_N78), .CK(clk), .Q(u5_prod1[78]) );
  DFF_X2 u5_prod_reg_78_ ( .D(u5_prod1[78]), .CK(clk), .Q(prod[78]), .QN(n4421) );
  DFF_X2 u5_prod1_reg_79_ ( .D(u5_N79), .CK(clk), .Q(u5_prod1[79]) );
  DFF_X2 u5_prod_reg_79_ ( .D(u5_prod1[79]), .CK(clk), .Q(prod[79]), .QN(n4436) );
  DFF_X2 u5_prod1_reg_80_ ( .D(u5_N80), .CK(clk), .Q(u5_prod1[80]) );
  DFF_X2 u5_prod_reg_80_ ( .D(u5_prod1[80]), .CK(clk), .Q(prod[80]), .QN(n4437) );
  DFF_X2 u5_prod1_reg_81_ ( .D(u5_N81), .CK(clk), .Q(u5_prod1[81]) );
  DFF_X2 u5_prod_reg_81_ ( .D(u5_prod1[81]), .CK(clk), .Q(prod[81]), .QN(n4427) );
  DFF_X2 u5_prod1_reg_82_ ( .D(u5_N82), .CK(clk), .Q(u5_prod1[82]) );
  DFF_X2 u5_prod_reg_82_ ( .D(u5_prod1[82]), .CK(clk), .Q(prod[82]), .QN(n4416) );
  DFF_X2 u5_prod1_reg_83_ ( .D(u5_N83), .CK(clk), .Q(u5_prod1[83]) );
  DFF_X2 u5_prod_reg_83_ ( .D(u5_prod1[83]), .CK(clk), .Q(prod[83]), .QN(n4420) );
  DFF_X2 u5_prod1_reg_84_ ( .D(u5_N84), .CK(clk), .Q(u5_prod1[84]) );
  DFF_X2 u5_prod_reg_84_ ( .D(u5_prod1[84]), .CK(clk), .QN(n4344) );
  DFF_X2 u5_prod1_reg_85_ ( .D(u5_N85), .CK(clk), .Q(u5_prod1[85]) );
  DFF_X2 u5_prod_reg_85_ ( .D(u5_prod1[85]), .CK(clk), .QN(n4404) );
  DFF_X2 u5_prod1_reg_86_ ( .D(u5_N86), .CK(clk), .Q(u5_prod1[86]) );
  DFF_X2 u5_prod_reg_86_ ( .D(u5_prod1[86]), .CK(clk), .QN(n4307) );
  DFF_X2 u5_prod1_reg_87_ ( .D(u5_N87), .CK(clk), .Q(u5_prod1[87]) );
  DFF_X2 u5_prod_reg_87_ ( .D(u5_prod1[87]), .CK(clk), .QN(n4294) );
  DFF_X2 u5_prod1_reg_88_ ( .D(u5_N88), .CK(clk), .Q(u5_prod1[88]) );
  DFF_X2 u5_prod_reg_88_ ( .D(u5_prod1[88]), .CK(clk), .Q(prod[88]), .QN(n4425) );
  DFF_X2 u5_prod1_reg_89_ ( .D(u5_N89), .CK(clk), .Q(u5_prod1[89]) );
  DFF_X2 u5_prod_reg_89_ ( .D(u5_prod1[89]), .CK(clk), .Q(prod[89]), .QN(n4411) );
  DFF_X2 u5_prod1_reg_90_ ( .D(u5_N90), .CK(clk), .Q(u5_prod1[90]) );
  DFF_X2 u5_prod_reg_90_ ( .D(u5_prod1[90]), .CK(clk), .QN(n4345) );
  DFF_X2 u5_prod1_reg_91_ ( .D(u5_N91), .CK(clk), .Q(u5_prod1[91]) );
  DFF_X2 u5_prod_reg_91_ ( .D(u5_prod1[91]), .CK(clk), .QN(n4405) );
  DFF_X2 u5_prod1_reg_92_ ( .D(u5_N92), .CK(clk), .Q(u5_prod1[92]) );
  DFF_X2 u5_prod_reg_92_ ( .D(u5_prod1[92]), .CK(clk), .QN(n4308) );
  DFF_X2 u5_prod1_reg_93_ ( .D(u5_N93), .CK(clk), .Q(u5_prod1[93]) );
  DFF_X2 u5_prod_reg_93_ ( .D(u5_prod1[93]), .CK(clk), .QN(n4295) );
  DFF_X2 u5_prod1_reg_94_ ( .D(u5_N94), .CK(clk), .Q(u5_prod1[94]) );
  DFF_X2 u5_prod_reg_94_ ( .D(u5_prod1[94]), .CK(clk), .Q(prod[94]), .QN(n4424) );
  DFF_X2 u5_prod1_reg_95_ ( .D(u5_N95), .CK(clk), .Q(u5_prod1[95]) );
  DFF_X2 u5_prod_reg_95_ ( .D(u5_prod1[95]), .CK(clk), .Q(prod[95]), .QN(n4408) );
  DFF_X2 u5_prod1_reg_96_ ( .D(u5_N96), .CK(clk), .Q(u5_prod1[96]) );
  DFF_X2 u5_prod_reg_96_ ( .D(u5_prod1[96]), .CK(clk), .Q(prod[96]), .QN(n4417) );
  DFF_X2 u5_prod1_reg_97_ ( .D(u5_N97), .CK(clk), .Q(u5_prod1[97]) );
  DFF_X2 u5_prod_reg_97_ ( .D(u5_prod1[97]), .CK(clk), .Q(prod[97]), .QN(n4431) );
  DFF_X2 u5_prod1_reg_98_ ( .D(u5_N98), .CK(clk), .Q(u5_prod1[98]) );
  DFF_X2 u5_prod_reg_98_ ( .D(u5_prod1[98]), .CK(clk), .Q(prod[98]), .QN(n4435) );
  DFF_X2 u5_prod1_reg_99_ ( .D(u5_N99), .CK(clk), .Q(u5_prod1[99]) );
  DFF_X2 u5_prod_reg_99_ ( .D(u5_prod1[99]), .CK(clk), .Q(prod[99]), .QN(n4433) );
  DFF_X2 u5_prod1_reg_100_ ( .D(u5_N100), .CK(clk), .Q(u5_prod1[100]) );
  DFF_X2 u5_prod_reg_100_ ( .D(u5_prod1[100]), .CK(clk), .Q(prod[100]), .QN(
        n4409) );
  DFF_X2 u5_prod1_reg_101_ ( .D(u5_N101), .CK(clk), .Q(u5_prod1[101]) );
  DFF_X2 u5_prod_reg_101_ ( .D(u5_prod1[101]), .CK(clk), .Q(prod[101]), .QN(
        n4418) );
  DFF_X2 u5_prod1_reg_102_ ( .D(u5_N102), .CK(clk), .Q(u5_prod1[102]) );
  DFF_X2 u5_prod_reg_102_ ( .D(u5_prod1[102]), .CK(clk), .QN(n4306) );
  DFF_X2 u5_prod1_reg_103_ ( .D(u5_N103), .CK(clk), .Q(u5_prod1[103]) );
  DFF_X2 u5_prod_reg_103_ ( .D(u5_prod1[103]), .CK(clk), .QN(n4403) );
  DFF_X2 u5_prod1_reg_104_ ( .D(u5_N104), .CK(clk), .Q(u5_prod1[104]) );
  DFF_X2 u5_prod_reg_104_ ( .D(u5_prod1[104]), .CK(clk), .QN(n4338) );
  DFF_X2 u5_prod1_reg_105_ ( .D(u5_N105), .CK(clk), .Q(u5_prod1[105]) );
  DFF_X2 u5_prod_reg_105_ ( .D(u5_prod1[105]), .CK(clk), .Q(prod[105]) );
  DFF_X2 u6_remainder_reg_0_ ( .D(u6_N0), .CK(clk), .Q(u6_remainder[0]) );
  DFF_X2 u6_rem_reg_0_ ( .D(u6_remainder[0]), .CK(clk), .Q(remainder[0]) );
  DFF_X2 u6_remainder_reg_1_ ( .D(u6_N1), .CK(clk), .Q(u6_remainder[1]) );
  DFF_X2 u6_rem_reg_1_ ( .D(u6_remainder[1]), .CK(clk), .Q(remainder[1]) );
  DFF_X2 u6_remainder_reg_2_ ( .D(u6_N2), .CK(clk), .Q(u6_remainder[2]) );
  DFF_X2 u6_rem_reg_2_ ( .D(u6_remainder[2]), .CK(clk), .Q(remainder[2]) );
  DFF_X2 u6_remainder_reg_3_ ( .D(u6_N3), .CK(clk), .Q(u6_remainder[3]) );
  DFF_X2 u6_rem_reg_3_ ( .D(u6_remainder[3]), .CK(clk), .Q(remainder[3]) );
  DFF_X2 u6_remainder_reg_4_ ( .D(u6_N4), .CK(clk), .Q(u6_remainder[4]) );
  DFF_X2 u6_rem_reg_4_ ( .D(u6_remainder[4]), .CK(clk), .Q(remainder[4]) );
  DFF_X2 u6_remainder_reg_5_ ( .D(u6_N5), .CK(clk), .Q(u6_remainder[5]) );
  DFF_X2 u6_rem_reg_5_ ( .D(u6_remainder[5]), .CK(clk), .Q(remainder[5]) );
  DFF_X2 u6_remainder_reg_6_ ( .D(u6_N6), .CK(clk), .Q(u6_remainder[6]) );
  DFF_X2 u6_rem_reg_6_ ( .D(u6_remainder[6]), .CK(clk), .Q(remainder[6]) );
  DFF_X2 u6_remainder_reg_7_ ( .D(u6_N7), .CK(clk), .Q(u6_remainder[7]) );
  DFF_X2 u6_rem_reg_7_ ( .D(u6_remainder[7]), .CK(clk), .Q(remainder[7]) );
  DFF_X2 u6_remainder_reg_8_ ( .D(u6_N8), .CK(clk), .Q(u6_remainder[8]) );
  DFF_X2 u6_rem_reg_8_ ( .D(u6_remainder[8]), .CK(clk), .Q(remainder[8]) );
  DFF_X2 u6_remainder_reg_9_ ( .D(u6_N9), .CK(clk), .Q(u6_remainder[9]) );
  DFF_X2 u6_rem_reg_9_ ( .D(u6_remainder[9]), .CK(clk), .Q(remainder[9]) );
  DFF_X2 u6_remainder_reg_10_ ( .D(u6_N10), .CK(clk), .Q(u6_remainder[10]) );
  DFF_X2 u6_rem_reg_10_ ( .D(u6_remainder[10]), .CK(clk), .Q(remainder[10]) );
  DFF_X2 u6_remainder_reg_11_ ( .D(u6_N11), .CK(clk), .Q(u6_remainder[11]) );
  DFF_X2 u6_rem_reg_11_ ( .D(u6_remainder[11]), .CK(clk), .Q(remainder[11]) );
  DFF_X2 u6_remainder_reg_12_ ( .D(u6_N12), .CK(clk), .Q(u6_remainder[12]) );
  DFF_X2 u6_rem_reg_12_ ( .D(u6_remainder[12]), .CK(clk), .Q(remainder[12]) );
  DFF_X2 u6_remainder_reg_13_ ( .D(u6_N13), .CK(clk), .Q(u6_remainder[13]) );
  DFF_X2 u6_rem_reg_13_ ( .D(u6_remainder[13]), .CK(clk), .Q(remainder[13]) );
  DFF_X2 u6_remainder_reg_14_ ( .D(u6_N14), .CK(clk), .Q(u6_remainder[14]) );
  DFF_X2 u6_rem_reg_14_ ( .D(u6_remainder[14]), .CK(clk), .Q(remainder[14]) );
  DFF_X2 u6_remainder_reg_15_ ( .D(u6_N15), .CK(clk), .Q(u6_remainder[15]) );
  DFF_X2 u6_rem_reg_15_ ( .D(u6_remainder[15]), .CK(clk), .Q(remainder[15]) );
  DFF_X2 u6_remainder_reg_16_ ( .D(u6_N16), .CK(clk), .Q(u6_remainder[16]) );
  DFF_X2 u6_rem_reg_16_ ( .D(u6_remainder[16]), .CK(clk), .Q(remainder[16]) );
  DFF_X2 u6_remainder_reg_17_ ( .D(u6_N17), .CK(clk), .Q(u6_remainder[17]) );
  DFF_X2 u6_rem_reg_17_ ( .D(u6_remainder[17]), .CK(clk), .Q(remainder[17]) );
  DFF_X2 u6_remainder_reg_18_ ( .D(u6_N18), .CK(clk), .Q(u6_remainder[18]) );
  DFF_X2 u6_rem_reg_18_ ( .D(u6_remainder[18]), .CK(clk), .Q(remainder[18]) );
  DFF_X2 u6_remainder_reg_19_ ( .D(u6_N19), .CK(clk), .Q(u6_remainder[19]) );
  DFF_X2 u6_rem_reg_19_ ( .D(u6_remainder[19]), .CK(clk), .Q(remainder[19]) );
  DFF_X2 u6_remainder_reg_20_ ( .D(u6_N20), .CK(clk), .Q(u6_remainder[20]) );
  DFF_X2 u6_rem_reg_20_ ( .D(u6_remainder[20]), .CK(clk), .Q(remainder[20]) );
  DFF_X2 u6_remainder_reg_21_ ( .D(u6_N21), .CK(clk), .Q(u6_remainder[21]) );
  DFF_X2 u6_rem_reg_21_ ( .D(u6_remainder[21]), .CK(clk), .Q(remainder[21]) );
  DFF_X2 u6_remainder_reg_22_ ( .D(u6_N22), .CK(clk), .Q(u6_remainder[22]) );
  DFF_X2 u6_rem_reg_22_ ( .D(u6_remainder[22]), .CK(clk), .Q(remainder[22]) );
  DFF_X2 u6_remainder_reg_23_ ( .D(u6_N23), .CK(clk), .Q(u6_remainder[23]) );
  DFF_X2 u6_rem_reg_23_ ( .D(u6_remainder[23]), .CK(clk), .Q(remainder[23]) );
  DFF_X2 u6_remainder_reg_24_ ( .D(u6_N24), .CK(clk), .Q(u6_remainder[24]) );
  DFF_X2 u6_rem_reg_24_ ( .D(u6_remainder[24]), .CK(clk), .Q(remainder[24]) );
  DFF_X2 u6_remainder_reg_25_ ( .D(u6_N25), .CK(clk), .Q(u6_remainder[25]) );
  DFF_X2 u6_rem_reg_25_ ( .D(u6_remainder[25]), .CK(clk), .Q(remainder[25]) );
  DFF_X2 u6_remainder_reg_26_ ( .D(u6_N26), .CK(clk), .Q(u6_remainder[26]) );
  DFF_X2 u6_rem_reg_26_ ( .D(u6_remainder[26]), .CK(clk), .Q(remainder[26]) );
  DFF_X2 u6_remainder_reg_27_ ( .D(u6_N27), .CK(clk), .Q(u6_remainder[27]) );
  DFF_X2 u6_rem_reg_27_ ( .D(u6_remainder[27]), .CK(clk), .Q(remainder[27]) );
  DFF_X2 u6_remainder_reg_28_ ( .D(u6_N28), .CK(clk), .Q(u6_remainder[28]) );
  DFF_X2 u6_rem_reg_28_ ( .D(u6_remainder[28]), .CK(clk), .Q(remainder[28]) );
  DFF_X2 u6_remainder_reg_29_ ( .D(u6_N29), .CK(clk), .Q(u6_remainder[29]) );
  DFF_X2 u6_rem_reg_29_ ( .D(u6_remainder[29]), .CK(clk), .Q(remainder[29]) );
  DFF_X2 u6_remainder_reg_30_ ( .D(u6_N30), .CK(clk), .Q(u6_remainder[30]) );
  DFF_X2 u6_rem_reg_30_ ( .D(u6_remainder[30]), .CK(clk), .Q(remainder[30]) );
  DFF_X2 u6_remainder_reg_31_ ( .D(u6_N31), .CK(clk), .Q(u6_remainder[31]) );
  DFF_X2 u6_rem_reg_31_ ( .D(u6_remainder[31]), .CK(clk), .Q(remainder[31]) );
  DFF_X2 u6_remainder_reg_32_ ( .D(u6_N32), .CK(clk), .Q(u6_remainder[32]) );
  DFF_X2 u6_rem_reg_32_ ( .D(u6_remainder[32]), .CK(clk), .Q(remainder[32]) );
  DFF_X2 u6_remainder_reg_33_ ( .D(u6_N33), .CK(clk), .Q(u6_remainder[33]) );
  DFF_X2 u6_rem_reg_33_ ( .D(u6_remainder[33]), .CK(clk), .Q(remainder[33]) );
  DFF_X2 u6_remainder_reg_34_ ( .D(u6_N34), .CK(clk), .Q(u6_remainder[34]) );
  DFF_X2 u6_rem_reg_34_ ( .D(u6_remainder[34]), .CK(clk), .Q(remainder[34]) );
  DFF_X2 u6_remainder_reg_35_ ( .D(u6_N35), .CK(clk), .Q(u6_remainder[35]) );
  DFF_X2 u6_rem_reg_35_ ( .D(u6_remainder[35]), .CK(clk), .Q(remainder[35]) );
  DFF_X2 u6_remainder_reg_36_ ( .D(u6_N36), .CK(clk), .Q(u6_remainder[36]) );
  DFF_X2 u6_rem_reg_36_ ( .D(u6_remainder[36]), .CK(clk), .Q(remainder[36]) );
  DFF_X2 u6_remainder_reg_37_ ( .D(u6_N37), .CK(clk), .Q(u6_remainder[37]) );
  DFF_X2 u6_rem_reg_37_ ( .D(u6_remainder[37]), .CK(clk), .Q(remainder[37]) );
  DFF_X2 u6_remainder_reg_38_ ( .D(u6_N38), .CK(clk), .Q(u6_remainder[38]) );
  DFF_X2 u6_rem_reg_38_ ( .D(u6_remainder[38]), .CK(clk), .Q(remainder[38]) );
  DFF_X2 u6_remainder_reg_39_ ( .D(u6_N39), .CK(clk), .Q(u6_remainder[39]) );
  DFF_X2 u6_rem_reg_39_ ( .D(u6_remainder[39]), .CK(clk), .Q(remainder[39]) );
  DFF_X2 u6_remainder_reg_40_ ( .D(u6_N40), .CK(clk), .Q(u6_remainder[40]) );
  DFF_X2 u6_rem_reg_40_ ( .D(u6_remainder[40]), .CK(clk), .Q(remainder[40]) );
  DFF_X2 u6_remainder_reg_41_ ( .D(u6_N41), .CK(clk), .Q(u6_remainder[41]) );
  DFF_X2 u6_rem_reg_41_ ( .D(u6_remainder[41]), .CK(clk), .Q(remainder[41]) );
  DFF_X2 u6_remainder_reg_42_ ( .D(u6_N42), .CK(clk), .Q(u6_remainder[42]) );
  DFF_X2 u6_rem_reg_42_ ( .D(u6_remainder[42]), .CK(clk), .Q(remainder[42]) );
  DFF_X2 u6_remainder_reg_43_ ( .D(u6_N43), .CK(clk), .Q(u6_remainder[43]) );
  DFF_X2 u6_rem_reg_43_ ( .D(u6_remainder[43]), .CK(clk), .Q(remainder[43]) );
  DFF_X2 u6_remainder_reg_44_ ( .D(u6_N44), .CK(clk), .Q(u6_remainder[44]) );
  DFF_X2 u6_rem_reg_44_ ( .D(u6_remainder[44]), .CK(clk), .Q(remainder[44]) );
  DFF_X2 u6_remainder_reg_45_ ( .D(u6_N45), .CK(clk), .Q(u6_remainder[45]) );
  DFF_X2 u6_rem_reg_45_ ( .D(u6_remainder[45]), .CK(clk), .Q(remainder[45]) );
  DFF_X2 u6_remainder_reg_46_ ( .D(u6_N46), .CK(clk), .Q(u6_remainder[46]) );
  DFF_X2 u6_rem_reg_46_ ( .D(u6_remainder[46]), .CK(clk), .Q(remainder[46]) );
  DFF_X2 u6_remainder_reg_47_ ( .D(u6_N47), .CK(clk), .Q(u6_remainder[47]) );
  DFF_X2 u6_rem_reg_47_ ( .D(u6_remainder[47]), .CK(clk), .Q(remainder[47]) );
  DFF_X2 u6_remainder_reg_48_ ( .D(u6_N48), .CK(clk), .Q(u6_remainder[48]) );
  DFF_X2 u6_rem_reg_48_ ( .D(u6_remainder[48]), .CK(clk), .Q(remainder[48]) );
  DFF_X2 u6_remainder_reg_49_ ( .D(u6_N49), .CK(clk), .Q(u6_remainder[49]) );
  DFF_X2 u6_rem_reg_49_ ( .D(u6_remainder[49]), .CK(clk), .Q(remainder[49]) );
  DFF_X2 u6_remainder_reg_50_ ( .D(u6_N50), .CK(clk), .Q(u6_remainder[50]) );
  DFF_X2 u6_rem_reg_50_ ( .D(u6_remainder[50]), .CK(clk), .Q(remainder[50]) );
  DFF_X2 u6_remainder_reg_51_ ( .D(u6_N51), .CK(clk), .Q(u6_remainder[51]) );
  DFF_X2 u6_rem_reg_51_ ( .D(u6_remainder[51]), .CK(clk), .Q(remainder[51]) );
  DFF_X2 u6_remainder_reg_52_ ( .D(u6_N52), .CK(clk), .Q(u6_remainder[52]) );
  DFF_X2 u6_rem_reg_52_ ( .D(u6_remainder[52]), .CK(clk), .Q(remainder[52]) );
  DFF_X2 u6_remainder_reg_55_ ( .D(u6_N55), .CK(clk), .Q(u6_remainder[55]) );
  DFF_X2 u6_rem_reg_55_ ( .D(u6_remainder[55]), .CK(clk), .Q(remainder[55]) );
  DFF_X2 u6_remainder_reg_56_ ( .D(u6_N56), .CK(clk), .Q(u6_remainder[56]) );
  DFF_X2 u6_rem_reg_56_ ( .D(u6_remainder[56]), .CK(clk), .Q(remainder[56]) );
  DFF_X2 u6_remainder_reg_57_ ( .D(u6_N57), .CK(clk), .Q(u6_remainder[57]) );
  DFF_X2 u6_rem_reg_57_ ( .D(u6_remainder[57]), .CK(clk), .Q(remainder[57]) );
  DFF_X2 u6_remainder_reg_58_ ( .D(u6_N58), .CK(clk), .Q(u6_remainder[58]) );
  DFF_X2 u6_rem_reg_58_ ( .D(u6_remainder[58]), .CK(clk), .Q(remainder[58]) );
  DFF_X2 u6_remainder_reg_59_ ( .D(u6_N59), .CK(clk), .Q(u6_remainder[59]) );
  DFF_X2 u6_rem_reg_59_ ( .D(u6_remainder[59]), .CK(clk), .Q(remainder[59]) );
  DFF_X2 u6_remainder_reg_60_ ( .D(u6_N60), .CK(clk), .Q(u6_remainder[60]) );
  DFF_X2 u6_rem_reg_60_ ( .D(u6_remainder[60]), .CK(clk), .Q(remainder[60]) );
  DFF_X2 u6_remainder_reg_61_ ( .D(u6_N61), .CK(clk), .Q(u6_remainder[61]) );
  DFF_X2 u6_rem_reg_61_ ( .D(u6_remainder[61]), .CK(clk), .Q(remainder[61]) );
  DFF_X2 u6_remainder_reg_62_ ( .D(u6_N62), .CK(clk), .Q(u6_remainder[62]) );
  DFF_X2 u6_rem_reg_62_ ( .D(u6_remainder[62]), .CK(clk), .Q(remainder[62]) );
  DFF_X2 u6_remainder_reg_63_ ( .D(u6_N63), .CK(clk), .Q(u6_remainder[63]) );
  DFF_X2 u6_rem_reg_63_ ( .D(u6_remainder[63]), .CK(clk), .Q(remainder[63]) );
  DFF_X2 u6_remainder_reg_64_ ( .D(u6_N64), .CK(clk), .Q(u6_remainder[64]) );
  DFF_X2 u6_rem_reg_64_ ( .D(u6_remainder[64]), .CK(clk), .Q(remainder[64]) );
  DFF_X2 u6_remainder_reg_65_ ( .D(u6_N65), .CK(clk), .Q(u6_remainder[65]) );
  DFF_X2 u6_rem_reg_65_ ( .D(u6_remainder[65]), .CK(clk), .Q(remainder[65]) );
  DFF_X2 u6_remainder_reg_66_ ( .D(u6_N66), .CK(clk), .Q(u6_remainder[66]) );
  DFF_X2 u6_rem_reg_66_ ( .D(u6_remainder[66]), .CK(clk), .Q(remainder[66]) );
  DFF_X2 u6_remainder_reg_67_ ( .D(u6_N67), .CK(clk), .Q(u6_remainder[67]) );
  DFF_X2 u6_rem_reg_67_ ( .D(u6_remainder[67]), .CK(clk), .Q(remainder[67]) );
  DFF_X2 u6_remainder_reg_68_ ( .D(u6_N68), .CK(clk), .Q(u6_remainder[68]) );
  DFF_X2 u6_rem_reg_68_ ( .D(u6_remainder[68]), .CK(clk), .Q(remainder[68]) );
  DFF_X2 u6_remainder_reg_69_ ( .D(u6_N69), .CK(clk), .Q(u6_remainder[69]) );
  DFF_X2 u6_rem_reg_69_ ( .D(u6_remainder[69]), .CK(clk), .Q(remainder[69]) );
  DFF_X2 u6_remainder_reg_70_ ( .D(u6_N70), .CK(clk), .Q(u6_remainder[70]) );
  DFF_X2 u6_rem_reg_70_ ( .D(u6_remainder[70]), .CK(clk), .Q(remainder[70]) );
  DFF_X2 u6_remainder_reg_71_ ( .D(u6_N71), .CK(clk), .Q(u6_remainder[71]) );
  DFF_X2 u6_rem_reg_71_ ( .D(u6_remainder[71]), .CK(clk), .Q(remainder[71]) );
  DFF_X2 u6_remainder_reg_72_ ( .D(u6_N72), .CK(clk), .Q(u6_remainder[72]) );
  DFF_X2 u6_rem_reg_72_ ( .D(u6_remainder[72]), .CK(clk), .Q(remainder[72]) );
  DFF_X2 u6_remainder_reg_73_ ( .D(u6_N73), .CK(clk), .Q(u6_remainder[73]) );
  DFF_X2 u6_rem_reg_73_ ( .D(u6_remainder[73]), .CK(clk), .Q(remainder[73]) );
  DFF_X2 u6_remainder_reg_74_ ( .D(u6_N74), .CK(clk), .Q(u6_remainder[74]) );
  DFF_X2 u6_rem_reg_74_ ( .D(u6_remainder[74]), .CK(clk), .Q(remainder[74]) );
  DFF_X2 u6_remainder_reg_75_ ( .D(u6_N75), .CK(clk), .Q(u6_remainder[75]) );
  DFF_X2 u6_rem_reg_75_ ( .D(u6_remainder[75]), .CK(clk), .Q(remainder[75]) );
  DFF_X2 u6_remainder_reg_76_ ( .D(u6_N76), .CK(clk), .Q(u6_remainder[76]) );
  DFF_X2 u6_rem_reg_76_ ( .D(u6_remainder[76]), .CK(clk), .Q(remainder[76]) );
  DFF_X2 u6_remainder_reg_77_ ( .D(u6_N77), .CK(clk), .Q(u6_remainder[77]) );
  DFF_X2 u6_rem_reg_77_ ( .D(u6_remainder[77]), .CK(clk), .Q(remainder[77]) );
  DFF_X2 u6_remainder_reg_78_ ( .D(u6_N78), .CK(clk), .Q(u6_remainder[78]) );
  DFF_X2 u6_rem_reg_78_ ( .D(u6_remainder[78]), .CK(clk), .Q(remainder[78]) );
  DFF_X2 u6_remainder_reg_79_ ( .D(u6_N79), .CK(clk), .Q(u6_remainder[79]) );
  DFF_X2 u6_rem_reg_79_ ( .D(u6_remainder[79]), .CK(clk), .Q(remainder[79]) );
  DFF_X2 u6_remainder_reg_80_ ( .D(u6_N80), .CK(clk), .Q(u6_remainder[80]) );
  DFF_X2 u6_rem_reg_80_ ( .D(u6_remainder[80]), .CK(clk), .Q(remainder[80]) );
  DFF_X2 u6_remainder_reg_81_ ( .D(u6_N81), .CK(clk), .Q(u6_remainder[81]) );
  DFF_X2 u6_rem_reg_81_ ( .D(u6_remainder[81]), .CK(clk), .Q(remainder[81]) );
  DFF_X2 u6_remainder_reg_82_ ( .D(u6_N82), .CK(clk), .Q(u6_remainder[82]) );
  DFF_X2 u6_rem_reg_82_ ( .D(u6_remainder[82]), .CK(clk), .Q(remainder[82]) );
  DFF_X2 u6_remainder_reg_83_ ( .D(u6_N83), .CK(clk), .Q(u6_remainder[83]) );
  DFF_X2 u6_rem_reg_83_ ( .D(u6_remainder[83]), .CK(clk), .Q(remainder[83]) );
  DFF_X2 u6_remainder_reg_84_ ( .D(u6_N84), .CK(clk), .Q(u6_remainder[84]) );
  DFF_X2 u6_rem_reg_84_ ( .D(u6_remainder[84]), .CK(clk), .Q(remainder[84]) );
  DFF_X2 u6_remainder_reg_85_ ( .D(u6_N85), .CK(clk), .Q(u6_remainder[85]) );
  DFF_X2 u6_rem_reg_85_ ( .D(u6_remainder[85]), .CK(clk), .Q(remainder[85]) );
  DFF_X2 u6_remainder_reg_86_ ( .D(u6_N86), .CK(clk), .Q(u6_remainder[86]) );
  DFF_X2 u6_rem_reg_86_ ( .D(u6_remainder[86]), .CK(clk), .Q(remainder[86]) );
  DFF_X2 u6_remainder_reg_87_ ( .D(u6_N87), .CK(clk), .Q(u6_remainder[87]) );
  DFF_X2 u6_rem_reg_87_ ( .D(u6_remainder[87]), .CK(clk), .Q(remainder[87]) );
  DFF_X2 u6_remainder_reg_88_ ( .D(u6_N88), .CK(clk), .Q(u6_remainder[88]) );
  DFF_X2 u6_rem_reg_88_ ( .D(u6_remainder[88]), .CK(clk), .Q(remainder[88]) );
  DFF_X2 u6_remainder_reg_89_ ( .D(u6_N89), .CK(clk), .Q(u6_remainder[89]) );
  DFF_X2 u6_rem_reg_89_ ( .D(u6_remainder[89]), .CK(clk), .Q(remainder[89]) );
  DFF_X2 u6_remainder_reg_90_ ( .D(u6_N90), .CK(clk), .Q(u6_remainder[90]) );
  DFF_X2 u6_rem_reg_90_ ( .D(u6_remainder[90]), .CK(clk), .Q(remainder[90]) );
  DFF_X2 u6_remainder_reg_91_ ( .D(u6_N91), .CK(clk), .Q(u6_remainder[91]) );
  DFF_X2 u6_rem_reg_91_ ( .D(u6_remainder[91]), .CK(clk), .Q(remainder[91]) );
  DFF_X2 u6_remainder_reg_92_ ( .D(u6_N92), .CK(clk), .Q(u6_remainder[92]) );
  DFF_X2 u6_rem_reg_92_ ( .D(u6_remainder[92]), .CK(clk), .Q(remainder[92]) );
  DFF_X2 u6_remainder_reg_93_ ( .D(u6_N93), .CK(clk), .Q(u6_remainder[93]) );
  DFF_X2 u6_rem_reg_93_ ( .D(u6_remainder[93]), .CK(clk), .Q(remainder[93]) );
  DFF_X2 u6_remainder_reg_94_ ( .D(u6_N94), .CK(clk), .Q(u6_remainder[94]) );
  DFF_X2 u6_rem_reg_94_ ( .D(u6_remainder[94]), .CK(clk), .Q(remainder[94]) );
  DFF_X2 u6_remainder_reg_95_ ( .D(u6_N95), .CK(clk), .Q(u6_remainder[95]) );
  DFF_X2 u6_rem_reg_95_ ( .D(u6_remainder[95]), .CK(clk), .Q(remainder[95]) );
  DFF_X2 u6_remainder_reg_96_ ( .D(u6_N96), .CK(clk), .Q(u6_remainder[96]) );
  DFF_X2 u6_rem_reg_96_ ( .D(u6_remainder[96]), .CK(clk), .Q(remainder[96]) );
  DFF_X2 u6_remainder_reg_97_ ( .D(u6_N97), .CK(clk), .Q(u6_remainder[97]) );
  DFF_X2 u6_rem_reg_97_ ( .D(u6_remainder[97]), .CK(clk), .Q(remainder[97]) );
  DFF_X2 u6_remainder_reg_98_ ( .D(u6_N98), .CK(clk), .Q(u6_remainder[98]) );
  DFF_X2 u6_rem_reg_98_ ( .D(u6_remainder[98]), .CK(clk), .Q(remainder[98]) );
  DFF_X2 u6_remainder_reg_99_ ( .D(u6_N99), .CK(clk), .Q(u6_remainder[99]) );
  DFF_X2 u6_rem_reg_99_ ( .D(u6_remainder[99]), .CK(clk), .Q(remainder[99]) );
  DFF_X2 u6_remainder_reg_100_ ( .D(u6_N100), .CK(clk), .Q(u6_remainder[100])
         );
  DFF_X2 u6_rem_reg_100_ ( .D(u6_remainder[100]), .CK(clk), .Q(remainder[100])
         );
  DFF_X2 u6_remainder_reg_101_ ( .D(u6_N101), .CK(clk), .Q(u6_remainder[101])
         );
  DFF_X2 u6_rem_reg_101_ ( .D(u6_remainder[101]), .CK(clk), .Q(remainder[101])
         );
  DFF_X2 u6_remainder_reg_102_ ( .D(u6_N102), .CK(clk), .Q(u6_remainder[102])
         );
  DFF_X2 u6_rem_reg_102_ ( .D(u6_remainder[102]), .CK(clk), .Q(remainder[102])
         );
  DFF_X2 u6_remainder_reg_103_ ( .D(u6_N103), .CK(clk), .Q(u6_remainder[103])
         );
  DFF_X2 u6_rem_reg_103_ ( .D(u6_remainder[103]), .CK(clk), .Q(remainder[103])
         );
  DFF_X2 u6_remainder_reg_104_ ( .D(u6_N104), .CK(clk), .Q(u6_remainder[104])
         );
  DFF_X2 u6_rem_reg_104_ ( .D(u6_remainder[104]), .CK(clk), .Q(remainder[104])
         );
  DFF_X2 u6_remainder_reg_105_ ( .D(u6_N105), .CK(clk), .Q(u6_remainder[105])
         );
  DFF_X2 u6_rem_reg_105_ ( .D(u6_remainder[105]), .CK(clk), .Q(remainder[105])
         );
  DFF_X2 u6_remainder_reg_106_ ( .D(u6_N106), .CK(clk), .Q(u6_remainder[106])
         );
  DFF_X2 u6_rem_reg_106_ ( .D(u6_remainder[106]), .CK(clk), .Q(remainder[106])
         );
  DFF_X2 u6_remainder_reg_107_ ( .D(u6_N107), .CK(clk), .Q(u6_remainder[107])
         );
  DFF_X2 u6_rem_reg_107_ ( .D(u6_remainder[107]), .CK(clk), .Q(remainder[107])
         );
  DFF_X2 u6_quo1_reg_0_ ( .D(u6_N0), .CK(clk), .Q(u6_quo1[0]) );
  DFF_X2 u6_quo_reg_0_ ( .D(u6_quo1[0]), .CK(clk), .Q(quo[0]) );
  DFF_X2 u6_quo1_reg_1_ ( .D(u6_N1), .CK(clk), .Q(u6_quo1[1]) );
  DFF_X2 u6_quo_reg_1_ ( .D(u6_quo1[1]), .CK(clk), .Q(quo[1]) );
  DFF_X2 u6_quo1_reg_2_ ( .D(u6_N2), .CK(clk), .Q(u6_quo1[2]) );
  DFF_X2 u6_quo_reg_2_ ( .D(u6_quo1[2]), .CK(clk), .Q(quo[2]) );
  DFF_X2 u6_quo1_reg_3_ ( .D(u6_N3), .CK(clk), .Q(u6_quo1[3]) );
  DFF_X2 u6_quo_reg_3_ ( .D(u6_quo1[3]), .CK(clk), .Q(quo[3]) );
  DFF_X2 u6_quo1_reg_4_ ( .D(u6_N4), .CK(clk), .Q(u6_quo1[4]) );
  DFF_X2 u6_quo_reg_4_ ( .D(u6_quo1[4]), .CK(clk), .Q(quo[4]) );
  DFF_X2 u6_quo1_reg_5_ ( .D(u6_N5), .CK(clk), .Q(u6_quo1[5]) );
  DFF_X2 u6_quo_reg_5_ ( .D(u6_quo1[5]), .CK(clk), .Q(quo[5]) );
  DFF_X2 u6_quo1_reg_6_ ( .D(u6_N6), .CK(clk), .Q(u6_quo1[6]) );
  DFF_X2 u6_quo_reg_6_ ( .D(u6_quo1[6]), .CK(clk), .Q(quo[6]) );
  DFF_X2 u6_quo1_reg_7_ ( .D(u6_N7), .CK(clk), .Q(u6_quo1[7]) );
  DFF_X2 u6_quo_reg_7_ ( .D(u6_quo1[7]), .CK(clk), .Q(quo[7]) );
  DFF_X2 u6_quo1_reg_8_ ( .D(u6_N8), .CK(clk), .Q(u6_quo1[8]) );
  DFF_X2 u6_quo_reg_8_ ( .D(u6_quo1[8]), .CK(clk), .Q(quo[8]) );
  DFF_X2 u6_quo1_reg_9_ ( .D(u6_N9), .CK(clk), .Q(u6_quo1[9]) );
  DFF_X2 u6_quo_reg_9_ ( .D(u6_quo1[9]), .CK(clk), .Q(quo[9]) );
  DFF_X2 u6_quo1_reg_10_ ( .D(u6_N10), .CK(clk), .Q(u6_quo1[10]) );
  DFF_X2 u6_quo_reg_10_ ( .D(u6_quo1[10]), .CK(clk), .Q(quo[10]) );
  DFF_X2 u6_quo1_reg_11_ ( .D(u6_N11), .CK(clk), .Q(u6_quo1[11]) );
  DFF_X2 u6_quo_reg_11_ ( .D(u6_quo1[11]), .CK(clk), .Q(quo[11]) );
  DFF_X2 u6_quo1_reg_12_ ( .D(u6_N12), .CK(clk), .Q(u6_quo1[12]) );
  DFF_X2 u6_quo_reg_12_ ( .D(u6_quo1[12]), .CK(clk), .Q(quo[12]) );
  DFF_X2 u6_quo1_reg_13_ ( .D(u6_N13), .CK(clk), .Q(u6_quo1[13]) );
  DFF_X2 u6_quo_reg_13_ ( .D(u6_quo1[13]), .CK(clk), .Q(quo[13]) );
  DFF_X2 u6_quo1_reg_14_ ( .D(u6_N14), .CK(clk), .Q(u6_quo1[14]) );
  DFF_X2 u6_quo_reg_14_ ( .D(u6_quo1[14]), .CK(clk), .Q(quo[14]) );
  DFF_X2 u6_quo1_reg_15_ ( .D(u6_N15), .CK(clk), .Q(u6_quo1[15]) );
  DFF_X2 u6_quo_reg_15_ ( .D(u6_quo1[15]), .CK(clk), .Q(quo[15]) );
  DFF_X2 u6_quo1_reg_16_ ( .D(u6_N16), .CK(clk), .Q(u6_quo1[16]) );
  DFF_X2 u6_quo_reg_16_ ( .D(u6_quo1[16]), .CK(clk), .Q(quo[16]) );
  DFF_X2 u6_quo1_reg_17_ ( .D(u6_N17), .CK(clk), .Q(u6_quo1[17]) );
  DFF_X2 u6_quo_reg_17_ ( .D(u6_quo1[17]), .CK(clk), .Q(quo[17]) );
  DFF_X2 u6_quo1_reg_18_ ( .D(u6_N18), .CK(clk), .Q(u6_quo1[18]) );
  DFF_X2 u6_quo_reg_18_ ( .D(u6_quo1[18]), .CK(clk), .Q(quo[18]) );
  DFF_X2 u6_quo1_reg_19_ ( .D(u6_N19), .CK(clk), .Q(u6_quo1[19]) );
  DFF_X2 u6_quo_reg_19_ ( .D(u6_quo1[19]), .CK(clk), .Q(quo[19]) );
  DFF_X2 u6_quo1_reg_20_ ( .D(u6_N20), .CK(clk), .Q(u6_quo1[20]) );
  DFF_X2 u6_quo_reg_20_ ( .D(u6_quo1[20]), .CK(clk), .Q(quo[20]) );
  DFF_X2 u6_quo1_reg_21_ ( .D(u6_N21), .CK(clk), .Q(u6_quo1[21]) );
  DFF_X2 u6_quo_reg_21_ ( .D(u6_quo1[21]), .CK(clk), .Q(quo[21]) );
  DFF_X2 u6_quo1_reg_22_ ( .D(u6_N22), .CK(clk), .Q(u6_quo1[22]) );
  DFF_X2 u6_quo_reg_22_ ( .D(u6_quo1[22]), .CK(clk), .Q(quo[22]) );
  DFF_X2 u6_quo1_reg_23_ ( .D(u6_N23), .CK(clk), .Q(u6_quo1[23]) );
  DFF_X2 u6_quo_reg_23_ ( .D(u6_quo1[23]), .CK(clk), .Q(quo[23]) );
  DFF_X2 u6_quo1_reg_24_ ( .D(u6_N24), .CK(clk), .Q(u6_quo1[24]) );
  DFF_X2 u6_quo_reg_24_ ( .D(u6_quo1[24]), .CK(clk), .Q(quo[24]) );
  DFF_X2 u6_quo1_reg_25_ ( .D(u6_N25), .CK(clk), .Q(u6_quo1[25]) );
  DFF_X2 u6_quo_reg_25_ ( .D(u6_quo1[25]), .CK(clk), .Q(quo[25]) );
  DFF_X2 u6_quo1_reg_26_ ( .D(u6_N26), .CK(clk), .Q(u6_quo1[26]) );
  DFF_X2 u6_quo_reg_26_ ( .D(u6_quo1[26]), .CK(clk), .Q(quo[26]) );
  DFF_X2 u6_quo1_reg_27_ ( .D(u6_N27), .CK(clk), .Q(u6_quo1[27]) );
  DFF_X2 u6_quo_reg_27_ ( .D(u6_quo1[27]), .CK(clk), .Q(quo[27]) );
  DFF_X2 u6_quo1_reg_28_ ( .D(u6_N28), .CK(clk), .Q(u6_quo1[28]) );
  DFF_X2 u6_quo_reg_28_ ( .D(u6_quo1[28]), .CK(clk), .Q(quo[28]) );
  DFF_X2 u6_quo1_reg_29_ ( .D(u6_N29), .CK(clk), .Q(u6_quo1[29]) );
  DFF_X2 u6_quo_reg_29_ ( .D(u6_quo1[29]), .CK(clk), .Q(quo[29]) );
  DFF_X2 u6_quo1_reg_30_ ( .D(u6_N30), .CK(clk), .Q(u6_quo1[30]) );
  DFF_X2 u6_quo_reg_30_ ( .D(u6_quo1[30]), .CK(clk), .Q(quo[30]) );
  DFF_X2 u6_quo1_reg_31_ ( .D(u6_N31), .CK(clk), .Q(u6_quo1[31]) );
  DFF_X2 u6_quo_reg_31_ ( .D(u6_quo1[31]), .CK(clk), .Q(quo[31]) );
  DFF_X2 u6_quo1_reg_32_ ( .D(u6_N32), .CK(clk), .Q(u6_quo1[32]) );
  DFF_X2 u6_quo_reg_32_ ( .D(u6_quo1[32]), .CK(clk), .Q(quo[32]) );
  DFF_X2 u6_quo1_reg_33_ ( .D(u6_N33), .CK(clk), .Q(u6_quo1[33]) );
  DFF_X2 u6_quo_reg_33_ ( .D(u6_quo1[33]), .CK(clk), .Q(quo[33]) );
  DFF_X2 u6_quo1_reg_34_ ( .D(u6_N34), .CK(clk), .Q(u6_quo1[34]) );
  DFF_X2 u6_quo_reg_34_ ( .D(u6_quo1[34]), .CK(clk), .Q(quo[34]) );
  DFF_X2 u6_quo1_reg_35_ ( .D(u6_N35), .CK(clk), .Q(u6_quo1[35]) );
  DFF_X2 u6_quo_reg_35_ ( .D(u6_quo1[35]), .CK(clk), .Q(quo[35]) );
  DFF_X2 u6_quo1_reg_36_ ( .D(u6_N36), .CK(clk), .Q(u6_quo1[36]) );
  DFF_X2 u6_quo_reg_36_ ( .D(u6_quo1[36]), .CK(clk), .Q(quo[36]) );
  DFF_X2 u6_quo1_reg_37_ ( .D(u6_N37), .CK(clk), .Q(u6_quo1[37]) );
  DFF_X2 u6_quo_reg_37_ ( .D(u6_quo1[37]), .CK(clk), .Q(quo[37]) );
  DFF_X2 u6_quo1_reg_38_ ( .D(u6_N38), .CK(clk), .Q(u6_quo1[38]) );
  DFF_X2 u6_quo_reg_38_ ( .D(u6_quo1[38]), .CK(clk), .Q(quo[38]) );
  DFF_X2 u6_quo1_reg_39_ ( .D(u6_N39), .CK(clk), .Q(u6_quo1[39]) );
  DFF_X2 u6_quo_reg_39_ ( .D(u6_quo1[39]), .CK(clk), .Q(quo[39]) );
  DFF_X2 u6_quo1_reg_40_ ( .D(u6_N40), .CK(clk), .Q(u6_quo1[40]) );
  DFF_X2 u6_quo_reg_40_ ( .D(u6_quo1[40]), .CK(clk), .Q(quo[40]) );
  DFF_X2 u6_quo1_reg_41_ ( .D(u6_N41), .CK(clk), .Q(u6_quo1[41]) );
  DFF_X2 u6_quo_reg_41_ ( .D(u6_quo1[41]), .CK(clk), .Q(quo[41]) );
  DFF_X2 u6_quo1_reg_42_ ( .D(u6_N42), .CK(clk), .Q(u6_quo1[42]) );
  DFF_X2 u6_quo_reg_42_ ( .D(u6_quo1[42]), .CK(clk), .Q(quo[42]) );
  DFF_X2 u6_quo1_reg_43_ ( .D(u6_N43), .CK(clk), .Q(u6_quo1[43]) );
  DFF_X2 u6_quo_reg_43_ ( .D(u6_quo1[43]), .CK(clk), .Q(quo[43]) );
  DFF_X2 u6_quo1_reg_44_ ( .D(u6_N44), .CK(clk), .Q(u6_quo1[44]) );
  DFF_X2 u6_quo_reg_44_ ( .D(u6_quo1[44]), .CK(clk), .Q(quo[44]) );
  DFF_X2 u6_quo1_reg_45_ ( .D(u6_N45), .CK(clk), .Q(u6_quo1[45]) );
  DFF_X2 u6_quo_reg_45_ ( .D(u6_quo1[45]), .CK(clk), .Q(quo[45]) );
  DFF_X2 u6_quo1_reg_46_ ( .D(u6_N46), .CK(clk), .Q(u6_quo1[46]) );
  DFF_X2 u6_quo_reg_46_ ( .D(u6_quo1[46]), .CK(clk), .Q(quo[46]) );
  DFF_X2 u6_quo1_reg_47_ ( .D(u6_N47), .CK(clk), .Q(u6_quo1[47]) );
  DFF_X2 u6_quo_reg_47_ ( .D(u6_quo1[47]), .CK(clk), .Q(quo[47]) );
  DFF_X2 u6_quo1_reg_48_ ( .D(u6_N48), .CK(clk), .Q(u6_quo1[48]) );
  DFF_X2 u6_quo_reg_48_ ( .D(u6_quo1[48]), .CK(clk), .Q(quo[48]) );
  DFF_X2 u6_quo1_reg_49_ ( .D(u6_N49), .CK(clk), .Q(u6_quo1[49]) );
  DFF_X2 u6_quo_reg_49_ ( .D(u6_quo1[49]), .CK(clk), .Q(quo[49]) );
  DFF_X2 u6_quo1_reg_50_ ( .D(u6_N50), .CK(clk), .Q(u6_quo1[50]) );
  DFF_X2 u6_quo_reg_50_ ( .D(u6_quo1[50]), .CK(clk), .Q(quo[50]) );
  DFF_X2 u6_quo1_reg_51_ ( .D(u6_N51), .CK(clk), .Q(u6_quo1[51]) );
  DFF_X2 u6_quo_reg_51_ ( .D(u6_quo1[51]), .CK(clk), .Q(quo[51]) );
  DFF_X2 u6_quo1_reg_52_ ( .D(u6_N52), .CK(clk), .Q(u6_quo1[52]) );
  DFF_X2 u6_quo_reg_52_ ( .D(u6_quo1[52]), .CK(clk), .Q(quo[52]) );
  DFF_X2 u6_quo1_reg_55_ ( .D(u6_N55), .CK(clk), .Q(u6_quo1[55]) );
  DFF_X2 u6_quo_reg_55_ ( .D(u6_quo1[55]), .CK(clk), .Q(quo[55]), .QN(n4398)
         );
  DFF_X2 u6_quo1_reg_56_ ( .D(u6_N56), .CK(clk), .Q(u6_quo1[56]) );
  DFF_X2 u6_quo_reg_56_ ( .D(u6_quo1[56]), .CK(clk), .Q(quo[56]) );
  DFF_X2 u6_quo1_reg_57_ ( .D(u6_N57), .CK(clk), .Q(u6_quo1[57]) );
  DFF_X2 u6_quo_reg_57_ ( .D(u6_quo1[57]), .CK(clk), .Q(quo[57]) );
  DFF_X2 u6_quo1_reg_58_ ( .D(u6_N58), .CK(clk), .Q(u6_quo1[58]) );
  DFF_X2 u6_quo_reg_58_ ( .D(u6_quo1[58]), .CK(clk), .Q(quo[58]) );
  DFF_X2 u6_quo1_reg_59_ ( .D(u6_N59), .CK(clk), .Q(u6_quo1[59]) );
  DFF_X2 u6_quo_reg_59_ ( .D(u6_quo1[59]), .CK(clk), .Q(quo[59]) );
  DFF_X2 u6_quo1_reg_60_ ( .D(u6_N60), .CK(clk), .Q(u6_quo1[60]) );
  DFF_X2 u6_quo_reg_60_ ( .D(u6_quo1[60]), .CK(clk), .Q(quo[60]) );
  DFF_X2 u6_quo1_reg_61_ ( .D(u6_N61), .CK(clk), .Q(u6_quo1[61]) );
  DFF_X2 u6_quo_reg_61_ ( .D(u6_quo1[61]), .CK(clk), .Q(quo[61]) );
  DFF_X2 u6_quo1_reg_62_ ( .D(u6_N62), .CK(clk), .Q(u6_quo1[62]) );
  DFF_X2 u6_quo_reg_62_ ( .D(u6_quo1[62]), .CK(clk), .Q(quo[62]) );
  DFF_X2 u6_quo1_reg_63_ ( .D(u6_N63), .CK(clk), .Q(u6_quo1[63]) );
  DFF_X2 u6_quo_reg_63_ ( .D(u6_quo1[63]), .CK(clk), .Q(quo[63]) );
  DFF_X2 u6_quo1_reg_64_ ( .D(u6_N64), .CK(clk), .Q(u6_quo1[64]) );
  DFF_X2 u6_quo_reg_64_ ( .D(u6_quo1[64]), .CK(clk), .Q(quo[64]) );
  DFF_X2 u6_quo1_reg_65_ ( .D(u6_N65), .CK(clk), .Q(u6_quo1[65]) );
  DFF_X2 u6_quo_reg_65_ ( .D(u6_quo1[65]), .CK(clk), .Q(quo[65]) );
  DFF_X2 u6_quo1_reg_66_ ( .D(u6_N66), .CK(clk), .Q(u6_quo1[66]) );
  DFF_X2 u6_quo_reg_66_ ( .D(u6_quo1[66]), .CK(clk), .Q(quo[66]) );
  DFF_X2 u6_quo1_reg_67_ ( .D(u6_N67), .CK(clk), .Q(u6_quo1[67]) );
  DFF_X2 u6_quo_reg_67_ ( .D(u6_quo1[67]), .CK(clk), .Q(quo[67]) );
  DFF_X2 u6_quo1_reg_68_ ( .D(u6_N68), .CK(clk), .Q(u6_quo1[68]) );
  DFF_X2 u6_quo_reg_68_ ( .D(u6_quo1[68]), .CK(clk), .Q(quo[68]) );
  DFF_X2 u6_quo1_reg_69_ ( .D(u6_N69), .CK(clk), .Q(u6_quo1[69]) );
  DFF_X2 u6_quo_reg_69_ ( .D(u6_quo1[69]), .CK(clk), .Q(quo[69]) );
  DFF_X2 u6_quo1_reg_70_ ( .D(u6_N70), .CK(clk), .Q(u6_quo1[70]) );
  DFF_X2 u6_quo_reg_70_ ( .D(u6_quo1[70]), .CK(clk), .Q(quo[70]) );
  DFF_X2 u6_quo1_reg_71_ ( .D(u6_N71), .CK(clk), .Q(u6_quo1[71]) );
  DFF_X2 u6_quo_reg_71_ ( .D(u6_quo1[71]), .CK(clk), .Q(quo[71]) );
  DFF_X2 u6_quo1_reg_72_ ( .D(u6_N72), .CK(clk), .Q(u6_quo1[72]) );
  DFF_X2 u6_quo_reg_72_ ( .D(u6_quo1[72]), .CK(clk), .Q(quo[72]) );
  DFF_X2 u6_quo1_reg_73_ ( .D(u6_N73), .CK(clk), .Q(u6_quo1[73]) );
  DFF_X2 u6_quo_reg_73_ ( .D(u6_quo1[73]), .CK(clk), .Q(quo[73]) );
  DFF_X2 u6_quo1_reg_74_ ( .D(u6_N74), .CK(clk), .Q(u6_quo1[74]) );
  DFF_X2 u6_quo_reg_74_ ( .D(u6_quo1[74]), .CK(clk), .Q(quo[74]) );
  DFF_X2 u6_quo1_reg_75_ ( .D(u6_N75), .CK(clk), .Q(u6_quo1[75]) );
  DFF_X2 u6_quo_reg_75_ ( .D(u6_quo1[75]), .CK(clk), .Q(quo[75]) );
  DFF_X2 u6_quo1_reg_76_ ( .D(u6_N76), .CK(clk), .Q(u6_quo1[76]) );
  DFF_X2 u6_quo_reg_76_ ( .D(u6_quo1[76]), .CK(clk), .Q(quo[76]) );
  DFF_X2 u6_quo1_reg_77_ ( .D(u6_N77), .CK(clk), .Q(u6_quo1[77]) );
  DFF_X2 u6_quo_reg_77_ ( .D(u6_quo1[77]), .CK(clk), .Q(quo[77]) );
  DFF_X2 u6_quo1_reg_78_ ( .D(u6_N78), .CK(clk), .Q(u6_quo1[78]) );
  DFF_X2 u6_quo_reg_78_ ( .D(u6_quo1[78]), .CK(clk), .Q(quo[78]) );
  DFF_X2 u6_quo1_reg_79_ ( .D(u6_N79), .CK(clk), .Q(u6_quo1[79]) );
  DFF_X2 u6_quo_reg_79_ ( .D(u6_quo1[79]), .CK(clk), .Q(quo[79]) );
  DFF_X2 u6_quo1_reg_80_ ( .D(u6_N80), .CK(clk), .Q(u6_quo1[80]) );
  DFF_X2 u6_quo_reg_80_ ( .D(u6_quo1[80]), .CK(clk), .Q(quo[80]) );
  DFF_X2 u6_quo1_reg_81_ ( .D(u6_N81), .CK(clk), .Q(u6_quo1[81]) );
  DFF_X2 u6_quo_reg_81_ ( .D(u6_quo1[81]), .CK(clk), .Q(quo[81]) );
  DFF_X2 u6_quo1_reg_82_ ( .D(u6_N82), .CK(clk), .Q(u6_quo1[82]) );
  DFF_X2 u6_quo_reg_82_ ( .D(u6_quo1[82]), .CK(clk), .Q(quo[82]) );
  DFF_X2 u6_quo1_reg_83_ ( .D(u6_N83), .CK(clk), .Q(u6_quo1[83]) );
  DFF_X2 u6_quo_reg_83_ ( .D(u6_quo1[83]), .CK(clk), .Q(quo[83]) );
  DFF_X2 u6_quo1_reg_84_ ( .D(u6_N84), .CK(clk), .Q(u6_quo1[84]) );
  DFF_X2 u6_quo_reg_84_ ( .D(u6_quo1[84]), .CK(clk), .Q(quo[84]) );
  DFF_X2 u6_quo1_reg_85_ ( .D(u6_N85), .CK(clk), .Q(u6_quo1[85]) );
  DFF_X2 u6_quo_reg_85_ ( .D(u6_quo1[85]), .CK(clk), .Q(quo[85]) );
  DFF_X2 u6_quo1_reg_86_ ( .D(u6_N86), .CK(clk), .Q(u6_quo1[86]) );
  DFF_X2 u6_quo_reg_86_ ( .D(u6_quo1[86]), .CK(clk), .Q(quo[86]) );
  DFF_X2 u6_quo1_reg_87_ ( .D(u6_N87), .CK(clk), .Q(u6_quo1[87]) );
  DFF_X2 u6_quo_reg_87_ ( .D(u6_quo1[87]), .CK(clk), .Q(quo[87]) );
  DFF_X2 u6_quo1_reg_88_ ( .D(u6_N88), .CK(clk), .Q(u6_quo1[88]) );
  DFF_X2 u6_quo_reg_88_ ( .D(u6_quo1[88]), .CK(clk), .Q(quo[88]) );
  DFF_X2 u6_quo1_reg_89_ ( .D(u6_N89), .CK(clk), .Q(u6_quo1[89]) );
  DFF_X2 u6_quo_reg_89_ ( .D(u6_quo1[89]), .CK(clk), .Q(quo[89]) );
  DFF_X2 u6_quo1_reg_90_ ( .D(u6_N90), .CK(clk), .Q(u6_quo1[90]) );
  DFF_X2 u6_quo_reg_90_ ( .D(u6_quo1[90]), .CK(clk), .Q(quo[90]) );
  DFF_X2 u6_quo1_reg_91_ ( .D(u6_N91), .CK(clk), .Q(u6_quo1[91]) );
  DFF_X2 u6_quo_reg_91_ ( .D(u6_quo1[91]), .CK(clk), .Q(quo[91]) );
  DFF_X2 u6_quo1_reg_92_ ( .D(u6_N92), .CK(clk), .Q(u6_quo1[92]) );
  DFF_X2 u6_quo_reg_92_ ( .D(u6_quo1[92]), .CK(clk), .Q(quo[92]) );
  DFF_X2 u6_quo1_reg_93_ ( .D(u6_N93), .CK(clk), .Q(u6_quo1[93]) );
  DFF_X2 u6_quo_reg_93_ ( .D(u6_quo1[93]), .CK(clk), .Q(quo[93]) );
  DFF_X2 u6_quo1_reg_94_ ( .D(u6_N94), .CK(clk), .Q(u6_quo1[94]) );
  DFF_X2 u6_quo_reg_94_ ( .D(u6_quo1[94]), .CK(clk), .Q(quo[94]) );
  DFF_X2 u6_quo1_reg_95_ ( .D(u6_N95), .CK(clk), .Q(u6_quo1[95]) );
  DFF_X2 u6_quo_reg_95_ ( .D(u6_quo1[95]), .CK(clk), .Q(quo[95]) );
  DFF_X2 u6_quo1_reg_96_ ( .D(u6_N96), .CK(clk), .Q(u6_quo1[96]) );
  DFF_X2 u6_quo_reg_96_ ( .D(u6_quo1[96]), .CK(clk), .Q(quo[96]) );
  DFF_X2 u6_quo1_reg_97_ ( .D(u6_N97), .CK(clk), .Q(u6_quo1[97]) );
  DFF_X2 u6_quo_reg_97_ ( .D(u6_quo1[97]), .CK(clk), .Q(quo[97]) );
  DFF_X2 u6_quo1_reg_98_ ( .D(u6_N98), .CK(clk), .Q(u6_quo1[98]) );
  DFF_X2 u6_quo_reg_98_ ( .D(u6_quo1[98]), .CK(clk), .Q(quo[98]) );
  DFF_X2 u6_quo1_reg_99_ ( .D(u6_N99), .CK(clk), .Q(u6_quo1[99]) );
  DFF_X2 u6_quo_reg_99_ ( .D(u6_quo1[99]), .CK(clk), .Q(quo[99]) );
  DFF_X2 u6_quo1_reg_100_ ( .D(u6_N100), .CK(clk), .Q(u6_quo1[100]) );
  DFF_X2 u6_quo_reg_100_ ( .D(u6_quo1[100]), .CK(clk), .Q(quo[100]) );
  DFF_X2 u6_quo1_reg_101_ ( .D(u6_N101), .CK(clk), .Q(u6_quo1[101]) );
  DFF_X2 u6_quo_reg_101_ ( .D(u6_quo1[101]), .CK(clk), .Q(quo[101]) );
  DFF_X2 u6_quo1_reg_102_ ( .D(u6_N102), .CK(clk), .Q(u6_quo1[102]) );
  DFF_X2 u6_quo_reg_102_ ( .D(u6_quo1[102]), .CK(clk), .Q(quo[102]) );
  DFF_X2 u6_quo1_reg_103_ ( .D(u6_N103), .CK(clk), .Q(u6_quo1[103]) );
  DFF_X2 u6_quo_reg_103_ ( .D(u6_quo1[103]), .CK(clk), .Q(quo[103]) );
  DFF_X2 u6_quo1_reg_104_ ( .D(u6_N104), .CK(clk), .Q(u6_quo1[104]) );
  DFF_X2 u6_quo_reg_104_ ( .D(u6_quo1[104]), .CK(clk), .Q(quo[104]) );
  DFF_X2 u6_quo1_reg_105_ ( .D(u6_N105), .CK(clk), .Q(u6_quo1[105]) );
  DFF_X2 u6_quo_reg_105_ ( .D(u6_quo1[105]), .CK(clk), .Q(quo[105]) );
  DFF_X2 u6_quo1_reg_106_ ( .D(u6_N106), .CK(clk), .Q(u6_quo1[106]) );
  DFF_X2 u6_quo_reg_106_ ( .D(u6_quo1[106]), .CK(clk), .Q(quo[106]) );
  DFF_X2 out_reg_55_ ( .D(N848), .CK(clk), .Q(out[55]) );
  DFF_X2 out_reg_56_ ( .D(N849), .CK(clk), .Q(out[56]) );
  DFF_X2 out_reg_54_ ( .D(N847), .CK(clk), .Q(out[54]) );
  DFF_X2 out_reg_57_ ( .D(N850), .CK(clk), .Q(out[57]) );
  DFF_X2 out_reg_59_ ( .D(N852), .CK(clk), .Q(out[59]) );
  DFF_X2 out_reg_58_ ( .D(N851), .CK(clk), .Q(out[58]) );
  DFF_X2 out_reg_53_ ( .D(N846), .CK(clk), .Q(out[53]) );
  DFF_X2 out_reg_52_ ( .D(N845), .CK(clk), .Q(out[52]) );
  DFF_X2 out_reg_62_ ( .D(N855), .CK(clk), .Q(out[62]) );
  DFF_X2 out_reg_61_ ( .D(N854), .CK(clk), .Q(out[61]) );
  DFF_X2 out_reg_60_ ( .D(N853), .CK(clk), .Q(out[60]) );
  DFF_X2 overflow_reg ( .D(N899), .CK(clk), .Q(overflow) );
  DFF_X2 out_reg_51_ ( .D(N844), .CK(clk), .Q(out[51]) );
  DFF_X2 out_reg_50_ ( .D(N843), .CK(clk), .Q(out[50]) );
  DFF_X2 out_reg_49_ ( .D(N842), .CK(clk), .Q(out[49]) );
  DFF_X2 out_reg_48_ ( .D(N841), .CK(clk), .Q(out[48]) );
  DFF_X2 out_reg_47_ ( .D(N840), .CK(clk), .Q(out[47]) );
  DFF_X2 out_reg_46_ ( .D(N839), .CK(clk), .Q(out[46]) );
  DFF_X2 out_reg_45_ ( .D(N838), .CK(clk), .Q(out[45]) );
  DFF_X2 out_reg_44_ ( .D(N837), .CK(clk), .Q(out[44]) );
  DFF_X2 out_reg_43_ ( .D(N836), .CK(clk), .Q(out[43]) );
  DFF_X2 out_reg_42_ ( .D(N835), .CK(clk), .Q(out[42]) );
  DFF_X2 out_reg_41_ ( .D(N834), .CK(clk), .Q(out[41]) );
  DFF_X2 out_reg_40_ ( .D(N833), .CK(clk), .Q(out[40]) );
  DFF_X2 out_reg_39_ ( .D(N832), .CK(clk), .Q(out[39]) );
  DFF_X2 out_reg_38_ ( .D(N831), .CK(clk), .Q(out[38]) );
  DFF_X2 out_reg_37_ ( .D(N830), .CK(clk), .Q(out[37]) );
  DFF_X2 out_reg_36_ ( .D(N829), .CK(clk), .Q(out[36]) );
  DFF_X2 out_reg_35_ ( .D(N828), .CK(clk), .Q(out[35]) );
  DFF_X2 out_reg_34_ ( .D(N827), .CK(clk), .Q(out[34]) );
  DFF_X2 out_reg_33_ ( .D(N826), .CK(clk), .Q(out[33]) );
  DFF_X2 out_reg_32_ ( .D(N825), .CK(clk), .Q(out[32]) );
  DFF_X2 out_reg_31_ ( .D(N824), .CK(clk), .Q(out[31]) );
  DFF_X2 out_reg_30_ ( .D(N823), .CK(clk), .Q(out[30]) );
  DFF_X2 out_reg_29_ ( .D(N822), .CK(clk), .Q(out[29]) );
  DFF_X2 out_reg_28_ ( .D(N821), .CK(clk), .Q(out[28]) );
  DFF_X2 out_reg_27_ ( .D(N820), .CK(clk), .Q(out[27]) );
  DFF_X2 out_reg_26_ ( .D(N819), .CK(clk), .Q(out[26]) );
  DFF_X2 out_reg_25_ ( .D(N818), .CK(clk), .Q(out[25]) );
  DFF_X2 out_reg_24_ ( .D(N817), .CK(clk), .Q(out[24]) );
  DFF_X2 out_reg_23_ ( .D(N816), .CK(clk), .Q(out[23]) );
  DFF_X2 out_reg_22_ ( .D(N815), .CK(clk), .Q(out[22]) );
  DFF_X2 out_reg_21_ ( .D(N814), .CK(clk), .Q(out[21]) );
  DFF_X2 out_reg_20_ ( .D(N813), .CK(clk), .Q(out[20]) );
  DFF_X2 out_reg_19_ ( .D(N812), .CK(clk), .Q(out[19]) );
  DFF_X2 out_reg_18_ ( .D(N811), .CK(clk), .Q(out[18]) );
  DFF_X2 out_reg_17_ ( .D(N810), .CK(clk), .Q(out[17]) );
  DFF_X2 out_reg_16_ ( .D(N809), .CK(clk), .Q(out[16]) );
  DFF_X2 out_reg_15_ ( .D(N808), .CK(clk), .Q(out[15]) );
  DFF_X2 out_reg_14_ ( .D(N807), .CK(clk), .Q(out[14]) );
  DFF_X2 out_reg_13_ ( .D(N806), .CK(clk), .Q(out[13]) );
  DFF_X2 out_reg_12_ ( .D(N805), .CK(clk), .Q(out[12]) );
  DFF_X2 out_reg_11_ ( .D(N804), .CK(clk), .Q(out[11]) );
  DFF_X2 out_reg_10_ ( .D(N803), .CK(clk), .Q(out[10]) );
  DFF_X2 out_reg_9_ ( .D(N802), .CK(clk), .Q(out[9]) );
  DFF_X2 out_reg_8_ ( .D(N801), .CK(clk), .Q(out[8]) );
  DFF_X2 out_reg_7_ ( .D(N800), .CK(clk), .Q(out[7]) );
  DFF_X2 out_reg_6_ ( .D(N799), .CK(clk), .Q(out[6]) );
  DFF_X2 out_reg_5_ ( .D(N798), .CK(clk), .Q(out[5]) );
  DFF_X2 out_reg_4_ ( .D(N797), .CK(clk), .Q(out[4]) );
  DFF_X2 out_reg_3_ ( .D(N796), .CK(clk), .Q(out[3]) );
  DFF_X2 out_reg_2_ ( .D(N795), .CK(clk), .Q(out[2]) );
  DFF_X2 out_reg_1_ ( .D(N794), .CK(clk), .Q(out[1]) );
  DFF_X2 inf_reg ( .D(N906), .CK(clk), .Q(inf) );
  DFF_X2 underflow_reg ( .D(N902), .CK(clk), .Q(underflow) );
  DFF_X2 ine_reg ( .D(N889), .CK(clk), .Q(ine) );
  DFF_X2 zero_reg ( .D(N911), .CK(clk), .Q(zero) );
  DFF_X2 out_reg_63_ ( .D(N875), .CK(clk), .Q(out[63]) );
  DFF_X2 out_reg_0_ ( .D(N793), .CK(clk), .Q(out[0]) );
  DFF_X2 u6_quo1_reg_107_ ( .D(u6_N107), .CK(clk), .Q(u6_quo1[107]) );
  DFF_X2 u6_quo_reg_107_ ( .D(u6_quo1[107]), .CK(clk), .Q(quo[107]) );
  FA_X1 u4_sub_412_U2_1 ( .A(div_opa_ldz_r2[1]), .B(n4314), .CI(
        u4_sub_412_carry[1]), .CO(u4_sub_412_carry[2]), .S(u4_div_shft4[1]) );
  FA_X1 u4_sub_412_U2_2 ( .A(div_opa_ldz_r2[2]), .B(n4438), .CI(
        u4_sub_412_carry[2]), .CO(u4_sub_412_carry[3]), .S(u4_div_shft4[2]) );
  FA_X1 u4_sub_412_U2_3 ( .A(div_opa_ldz_r2[3]), .B(n4316), .CI(
        u4_sub_412_carry[3]), .CO(u4_sub_412_carry[4]), .S(u4_div_shft4[3]) );
  FA_X1 u4_sub_412_U2_4 ( .A(div_opa_ldz_r2[4]), .B(n4299), .CI(
        u4_sub_412_carry[4]), .CO(u4_sub_412_carry[5]), .S(u4_div_shft4[4]) );
  FA_X1 u4_add_411_U1_1 ( .A(div_opa_ldz_r2[1]), .B(exp_r[1]), .CI(
        u4_add_411_carry[1]), .CO(u4_add_411_carry[2]), .S(u4_div_shft3_1_) );
  FA_X1 u4_add_411_U1_2 ( .A(div_opa_ldz_r2[2]), .B(n4315), .CI(
        u4_add_411_carry[2]), .CO(u4_add_411_carry[3]), .S(u4_div_shft3_2_) );
  FA_X1 u4_add_411_U1_3 ( .A(div_opa_ldz_r2[3]), .B(n4655), .CI(
        u4_add_411_carry[3]), .CO(u4_add_411_carry[4]), .S(u4_div_shft3_3_) );
  FA_X1 u4_add_411_U1_4 ( .A(div_opa_ldz_r2[4]), .B(n4282), .CI(
        u4_add_411_carry[4]), .CO(u4_add_411_carry[5]), .S(u4_div_shft3_4_) );
  FA_X1 u4_sub_409_U2_1 ( .A(exp_r[1]), .B(n4446), .CI(u4_sub_409_carry[1]), 
        .CO(u4_sub_409_carry[2]), .S(u4_div_scht1a[1]) );
  FA_X1 u4_sub_409_U2_2 ( .A(n4315), .B(n4444), .CI(u4_sub_409_carry[2]), .CO(
        u4_sub_409_carry[3]), .S(u4_div_scht1a[2]) );
  FA_X1 u4_sub_409_U2_3 ( .A(n4655), .B(n4443), .CI(u4_sub_409_carry[3]), .CO(
        u4_sub_409_carry[4]), .S(u4_div_scht1a[3]) );
  FA_X1 u4_sub_409_U2_4 ( .A(n4282), .B(n4445), .CI(u4_sub_409_carry[4]), .CO(
        u4_sub_409_carry[5]), .S(u4_div_scht1a[4]) );
  FA_X1 sub_1_root_sub_0_root_u4_add_497_U2_1 ( .A(exp_r[1]), .B(n4446), .CI(
        sub_1_root_sub_0_root_u4_add_497_carry[1]), .CO(
        sub_1_root_sub_0_root_u4_add_497_carry[2]), .S(u4_ldz_dif_1_) );
  FA_X1 sub_1_root_sub_0_root_u4_add_497_U2_2 ( .A(n4315), .B(n4444), .CI(
        sub_1_root_sub_0_root_u4_add_497_carry[2]), .CO(
        sub_1_root_sub_0_root_u4_add_497_carry[3]), .S(u4_ldz_dif_2_) );
  FA_X1 sub_1_root_sub_0_root_u4_add_497_U2_3 ( .A(n4655), .B(n4443), .CI(
        sub_1_root_sub_0_root_u4_add_497_carry[3]), .CO(
        sub_1_root_sub_0_root_u4_add_497_carry[4]), .S(u4_ldz_dif_3_) );
  FA_X1 sub_1_root_sub_0_root_u4_add_497_U2_4 ( .A(n4282), .B(n4445), .CI(
        sub_1_root_sub_0_root_u4_add_497_carry[4]), .CO(
        sub_1_root_sub_0_root_u4_add_497_carry[5]), .S(u4_ldz_dif_4_) );
  NAND2_X2 U3379 ( .A1(quo[2]), .A2(n4563), .ZN(n4027) );
  NAND2_X2 U3380 ( .A1(quo[106]), .A2(n4575), .ZN(n4111) );
  NAND2_X2 U3381 ( .A1(quo[1]), .A2(n4563), .ZN(n3977) );
  NAND2_X2 U3382 ( .A1(quo[105]), .A2(n4574), .ZN(n4113) );
  NOR2_X4 U3383 ( .A1(remainder[56]), .A2(remainder[55]), .ZN(n4152) );
  NOR2_X4 U3384 ( .A1(remainder[51]), .A2(remainder[52]), .ZN(n4151) );
  NOR3_X2 U3385 ( .A1(n3741), .A2(n3849), .A3(n3551), .ZN(n3803) );
  NAND3_X2 U3386 ( .A1(n3851), .A2(n3834), .A3(rmode_r3[1]), .ZN(n3850) );
  NAND3_X2 U3387 ( .A1(n3557), .A2(n2434), .A3(sign), .ZN(n3851) );
  AOI222_X1 U3388 ( .A1(n4600), .A2(n2483), .B1(n4349), .B2(n6342), .C1(
        div_opa_ldz_r2[0]), .C2(n2498), .ZN(n2513) );
  AOI222_X1 U3389 ( .A1(u4_fi_ldz_1_), .A2(n2489), .B1(exp_r[1]), .B2(n2483), 
        .C1(u4_div_scht1a[1]), .C2(n2484), .ZN(n2503) );
  OAI21_X2 U3390 ( .B1(n3767), .B2(n4355), .A(n3768), .ZN(n3477) );
  AOI21_X2 U3391 ( .B1(n6305), .B2(n3773), .A(n3774), .ZN(n3767) );
  NOR3_X2 U3392 ( .A1(n2465), .A2(n2459), .A3(n2462), .ZN(n3856) );
  NAND3_X2 U3393 ( .A1(u4_exp_out_0_), .A2(u4_exp_out_10_), .A3(u4_exp_out_9_), 
        .ZN(n3858) );
  NOR3_X2 U3394 ( .A1(fract_denorm[93]), .A2(fract_denorm[94]), .A3(n6357), 
        .ZN(n2707) );
  AOI21_X2 U3395 ( .B1(n2434), .B2(n3557), .A(n3849), .ZN(n3852) );
  NOR3_X2 U3396 ( .A1(n2514), .A2(n2515), .A3(n4355), .ZN(n2498) );
  NAND3_X2 U3397 ( .A1(n2709), .A2(n6413), .A3(n2555), .ZN(n2602) );
  NOR3_X2 U3398 ( .A1(fract_denorm[83]), .A2(fract_denorm[84]), .A3(n6375), 
        .ZN(n2644) );
  AOI21_X2 U3399 ( .B1(n2700), .B2(n6347), .A(n2701), .ZN(n2699) );
  NAND3_X2 U3400 ( .A1(n2660), .A2(n6422), .A3(n2600), .ZN(n2615) );
  NOR3_X2 U3401 ( .A1(fract_denorm[96]), .A2(fract_denorm[97]), .A3(
        fract_denorm[95]), .ZN(n2738) );
  NOR3_X2 U3402 ( .A1(n2635), .A2(n6442), .A3(n6329), .ZN(n2555) );
  AOI21_X2 U3403 ( .B1(n6466), .B2(exp_ovf_r[0]), .A(n5912), .ZN(n3777) );
  AOI21_X2 U3404 ( .B1(u4_N6251), .B2(n3557), .A(n5912), .ZN(n3776) );
  AOI222_X1 U3405 ( .A1(n3829), .A2(u4_exp_out_10_), .B1(n3802), .B2(
        u4_exp_next_mi_10_), .C1(u4_exp_out_pl1_10_), .C2(n3805), .ZN(n3842)
         );
  AOI222_X1 U3406 ( .A1(n3829), .A2(u4_exp_out_0_), .B1(n3802), .B2(
        u4_exp_next_mi_0_), .C1(u4_exp_out_pl1_0_), .C2(n3805), .ZN(n3828) );
  AOI211_X2 U3407 ( .C1(n4452), .C2(n3476), .A(n2480), .B(u4_exp_in_mi1_11_), 
        .ZN(n2506) );
  NAND3_X2 U3408 ( .A1(n4452), .A2(n3489), .A3(n6447), .ZN(n2518) );
  NOR3_X2 U3409 ( .A1(n6393), .A2(fract_denorm[66]), .A3(n6335), .ZN(n2562) );
  NAND3_X2 U3410 ( .A1(n2609), .A2(n2585), .A3(n2710), .ZN(n2641) );
  NOR3_X2 U3411 ( .A1(n2634), .A2(n6440), .A3(n2632), .ZN(n2639) );
  NOR3_X2 U3412 ( .A1(n2635), .A2(n2636), .A3(n6329), .ZN(n2611) );
  NOR3_X2 U3413 ( .A1(n2648), .A2(n2649), .A3(n2650), .ZN(n2626) );
  NOR3_X2 U3414 ( .A1(fract_denorm[103]), .A2(fract_denorm[104]), .A3(n2662), 
        .ZN(n2761) );
  OAI21_X2 U3415 ( .B1(n4540), .B2(n3787), .A(n3788), .ZN(n3786) );
  OAI21_X2 U3416 ( .B1(n3789), .B2(n3783), .A(n3790), .ZN(n3785) );
  NOR3_X2 U3417 ( .A1(n2515), .A2(n6465), .A3(n4355), .ZN(n2484) );
  AOI211_X2 U3418 ( .C1(n2686), .C2(n4653), .A(n2687), .B(n2688), .ZN(n2673)
         );
  OAI21_X2 U3419 ( .B1(fract_denorm[105]), .B2(n6096), .A(n2514), .ZN(n3963)
         );
  NOR3_X2 U3420 ( .A1(n3608), .A2(n3609), .A3(n3610), .ZN(n3570) );
  NOR2_X2 U3421 ( .A1(n2434), .A2(n3304), .ZN(n3302) );
  NAND3_X2 U3422 ( .A1(n3456), .A2(n3461), .A3(n3342), .ZN(n3463) );
  AOI21_X2 U3423 ( .B1(n6305), .B2(n6459), .A(n3463), .ZN(n3465) );
  OAI21_X2 U3424 ( .B1(n3318), .B2(n3319), .A(n3320), .ZN(n3316) );
  OAI21_X2 U3425 ( .B1(n3551), .B2(n6094), .A(n3552), .ZN(n3550) );
  NOR3_X2 U3426 ( .A1(n3555), .A2(n3556), .A3(n3477), .ZN(n3553) );
  AOI222_X1 U3427 ( .A1(n2679), .A2(fract_denorm[57]), .B1(n2600), .B2(n6424), 
        .C1(n6327), .C2(n6438), .ZN(n2714) );
  NOR3_X2 U3428 ( .A1(n2690), .A2(n2691), .A3(n2664), .ZN(n2712) );
  AOI211_X2 U3429 ( .C1(n2716), .C2(n6362), .A(n4652), .B(n2717), .ZN(n2715)
         );
  NOR2_X2 U3430 ( .A1(n6362), .A2(n2399), .ZN(n2391) );
  NOR2_X2 U3431 ( .A1(n2399), .A2(n6094), .ZN(n2401) );
  INV_X4 U3432 ( .A(n4619), .ZN(n4608) );
  NOR3_X2 U3433 ( .A1(n6440), .A2(n6445), .A3(n6346), .ZN(n3872) );
  AOI21_X2 U3434 ( .B1(n3495), .B2(n4540), .A(n3544), .ZN(n3882) );
  NOR3_X2 U3435 ( .A1(exp_r[1]), .A2(n4655), .A3(n4315), .ZN(n3907) );
  INV_X4 U3436 ( .A(n4616), .ZN(n4613) );
  INV_X4 U3437 ( .A(n4627), .ZN(n4625) );
  INV_X4 U3438 ( .A(n4619), .ZN(n4609) );
  INV_X4 U3439 ( .A(n4627), .ZN(n4624) );
  INV_X4 U3440 ( .A(n4616), .ZN(n4614) );
  NAND2_X2 U3441 ( .A1(n4603), .A2(n6303), .ZN(n3052) );
  NOR2_X2 U3442 ( .A1(n2955), .A2(n6238), .ZN(n2977) );
  NAND3_X2 U3443 ( .A1(n3037), .A2(n3038), .A3(n3039), .ZN(n3036) );
  NAND3_X2 U3444 ( .A1(n3041), .A2(n3042), .A3(n3043), .ZN(n3040) );
  NAND3_X2 U3445 ( .A1(n3045), .A2(n3046), .A3(n3047), .ZN(n3044) );
  NOR2_X2 U3446 ( .A1(u1_exp_lt_27), .A2(u1_exp_diff_4_), .ZN(n3012) );
  NOR2_X2 U3447 ( .A1(n2954), .A2(u1_adj_op_51_), .ZN(n2976) );
  NOR2_X2 U3448 ( .A1(u1_exp_lt_27), .A2(u1_exp_diff_3_), .ZN(n3001) );
  NOR2_X2 U3449 ( .A1(n3004), .A2(n6225), .ZN(n3002) );
  NOR3_X2 U3450 ( .A1(n3004), .A2(n6224), .A3(n3012), .ZN(n3011) );
  NOR3_X2 U3451 ( .A1(fract_denorm[77]), .A2(fract_denorm[78]), .A3(n6385), 
        .ZN(n2728) );
  NAND3_X2 U3452 ( .A1(n6353), .A2(n6354), .A3(n2707), .ZN(n2599) );
  NOR3_X2 U3453 ( .A1(n6409), .A2(n6367), .A3(n6410), .ZN(n2668) );
  NOR3_X2 U3454 ( .A1(n6344), .A2(n6345), .A3(n6441), .ZN(n3878) );
  NOR3_X2 U3455 ( .A1(n3869), .A2(n3870), .A3(n3871), .ZN(n3868) );
  NAND3_X2 U3456 ( .A1(n2683), .A2(n2718), .A3(n2767), .ZN(n3870) );
  NAND3_X2 U3457 ( .A1(n3171), .A2(n2751), .A3(n6400), .ZN(n3871) );
  OAI21_X2 U3458 ( .B1(n3882), .B2(n3883), .A(n3884), .ZN(n3880) );
  NOR3_X2 U3459 ( .A1(n3906), .A2(n3771), .A3(n4540), .ZN(n3883) );
  NAND3_X2 U3460 ( .A1(n3885), .A2(n6337), .A3(exp_ovf_r[1]), .ZN(n3884) );
  NOR3_X2 U3461 ( .A1(n6416), .A2(n6417), .A3(n6418), .ZN(n2670) );
  NOR3_X2 U3462 ( .A1(fract_denorm[53]), .A2(fract_denorm[54]), .A3(n6372), 
        .ZN(n2698) );
  NOR3_X2 U3463 ( .A1(n6380), .A2(n2592), .A3(n6393), .ZN(n4016) );
  NOR3_X2 U3464 ( .A1(fract_denorm[75]), .A2(fract_denorm[76]), .A3(n6382), 
        .ZN(n2560) );
  NOR3_X2 U3465 ( .A1(u4_N6040), .A2(u4_N6042), .A3(u4_N6041), .ZN(n3948) );
  NOR3_X2 U3466 ( .A1(u4_N6043), .A2(u4_N6045), .A3(u4_N6044), .ZN(n3949) );
  NOR3_X2 U3467 ( .A1(u4_N6046), .A2(u4_N6048), .A3(u4_N6047), .ZN(n3950) );
  NOR3_X2 U3468 ( .A1(u4_N6053), .A2(u4_N6055), .A3(u4_N6054), .ZN(n3952) );
  NOR3_X2 U3469 ( .A1(u4_N6060), .A2(u4_N6062), .A3(u4_N6061), .ZN(n3954) );
  NOR3_X2 U3470 ( .A1(u4_N6027), .A2(u4_N6029), .A3(u4_N6028), .ZN(n3944) );
  NOR3_X2 U3471 ( .A1(u4_N6030), .A2(u4_N6032), .A3(u4_N6031), .ZN(n3945) );
  NOR3_X2 U3472 ( .A1(u4_N6033), .A2(u4_N6035), .A3(u4_N6034), .ZN(n3946) );
  NOR3_X2 U3473 ( .A1(u4_N6014), .A2(u4_N6016), .A3(u4_N6015), .ZN(n3940) );
  NOR3_X2 U3474 ( .A1(u4_N6017), .A2(u4_N6019), .A3(u4_N6018), .ZN(n3941) );
  NOR3_X2 U3475 ( .A1(u4_N6020), .A2(u4_N6022), .A3(u4_N6021), .ZN(n3942) );
  NAND3_X2 U3476 ( .A1(n2410), .A2(n2406), .A3(n2413), .ZN(n3505) );
  NOR3_X2 U3477 ( .A1(u4_fract_out_12_), .A2(u4_fract_out_14_), .A3(
        u4_fract_out_13_), .ZN(n3902) );
  NOR3_X2 U3478 ( .A1(u4_fract_out_36_), .A2(u4_fract_out_38_), .A3(
        u4_fract_out_37_), .ZN(n3892) );
  NOR3_X2 U3479 ( .A1(u4_fract_out_48_), .A2(u4_fract_out_4_), .A3(
        u4_fract_out_49_), .ZN(n3896) );
  NOR3_X2 U3480 ( .A1(u4_fract_out_24_), .A2(u4_fract_out_26_), .A3(
        u4_fract_out_25_), .ZN(n3904) );
  OAI21_X2 U3481 ( .B1(u4_fract_out_0_), .B2(n3853), .A(n3854), .ZN(n3743) );
  AOI21_X2 U3482 ( .B1(sign), .B2(rmode_r3[1]), .A(n6305), .ZN(n3736) );
  NOR3_X2 U3483 ( .A1(n4789), .A2(u4_fi_ldz_2a_6_), .A3(u4_fi_ldz_2a_5_), .ZN(
        u4_N6251) );
  NOR2_X2 U3484 ( .A1(n2434), .A2(n6307), .ZN(n3737) );
  NAND3_X2 U3485 ( .A1(n6305), .A2(n4540), .A3(n3849), .ZN(n3855) );
  AOI222_X1 U3486 ( .A1(n4540), .A2(opb_inf), .B1(n3297), .B2(opa_00), .C1(
        n6316), .C2(opb_00), .ZN(n3745) );
  NOR2_X2 U3487 ( .A1(u1_exp_lt_27), .A2(u1_exp_diff_5_), .ZN(n3004) );
  INV_X4 U3488 ( .A(n4604), .ZN(n4632) );
  INV_X4 U3489 ( .A(n4605), .ZN(n4604) );
  INV_X4 U3490 ( .A(u1_expa_lt_expb), .ZN(n4605) );
  AOI222_X1 U3491 ( .A1(n6213), .A2(n2971), .B1(n6212), .B2(n2972), .C1(n6219), 
        .C2(n2973), .ZN(n2970) );
  NOR2_X2 U3492 ( .A1(n2991), .A2(u1_adj_op_42_), .ZN(n2959) );
  NOR2_X2 U3493 ( .A1(n2992), .A2(u1_adj_op_38_), .ZN(n2957) );
  NAND3_X2 U3494 ( .A1(n6224), .A2(n3003), .A3(n3002), .ZN(n2958) );
  NOR2_X2 U3495 ( .A1(n2971), .A2(u1_adj_op_28_), .ZN(n2996) );
  NAND3_X2 U3496 ( .A1(n6217), .A2(n6224), .A3(n3002), .ZN(n2960) );
  AOI21_X2 U3497 ( .B1(n2976), .B2(n6273), .A(n3001), .ZN(n3008) );
  NOR3_X2 U3498 ( .A1(n3012), .A2(n6217), .A3(n3004), .ZN(n3009) );
  NOR2_X2 U3499 ( .A1(n2978), .A2(u1_adj_op_44_), .ZN(n3005) );
  NOR2_X2 U3500 ( .A1(n2979), .A2(n6243), .ZN(n3006) );
  NOR2_X2 U3501 ( .A1(n3010), .A2(n6236), .ZN(n2988) );
  NOR2_X2 U3502 ( .A1(n3000), .A2(n6247), .ZN(n2986) );
  NAND3_X2 U3503 ( .A1(n6217), .A2(n3001), .A3(n3002), .ZN(n2968) );
  NAND3_X2 U3504 ( .A1(n3003), .A2(n3001), .A3(n3002), .ZN(n2966) );
  AOI222_X1 U3505 ( .A1(n4655), .A2(n2483), .B1(u4_f2i_shft_3_), .B2(n6342), 
        .C1(div_opa_ldz_r2[3]), .C2(n2498), .ZN(n2500) );
  NOR2_X2 U3506 ( .A1(n6465), .A2(u4_exp_in_pl1_1_), .ZN(n2510) );
  AOI222_X1 U3507 ( .A1(n4315), .A2(n2483), .B1(u4_f2i_shft_2_), .B2(n6342), 
        .C1(div_opa_ldz_r2[2]), .C2(n2498), .ZN(n2502) );
  AOI222_X1 U3508 ( .A1(n4282), .A2(n2483), .B1(u4_f2i_shft_4_), .B2(n6342), 
        .C1(div_opa_ldz_r2[4]), .C2(n2498), .ZN(n2497) );
  AOI222_X1 U3509 ( .A1(u4_div_scht1a[5]), .A2(n2484), .B1(u4_f2i_shft_5_), 
        .B2(n6342), .C1(n4290), .C2(n2483), .ZN(n2494) );
  NAND3_X2 U3510 ( .A1(n3173), .A2(n2729), .A3(n2706), .ZN(n2771) );
  AOI21_X2 U3511 ( .B1(n6371), .B2(n6373), .A(n6326), .ZN(n2591) );
  NOR3_X2 U3512 ( .A1(n6334), .A2(n6401), .A3(n2592), .ZN(n2590) );
  NOR3_X2 U3513 ( .A1(fract_denorm[64]), .A2(fract_denorm[65]), .A3(
        fract_denorm[63]), .ZN(n2735) );
  NOR3_X2 U3514 ( .A1(fract_denorm[61]), .A2(fract_denorm[62]), .A3(n6391), 
        .ZN(n2705) );
  NAND3_X2 U3515 ( .A1(n2560), .A2(fract_denorm[74]), .A3(n6325), .ZN(n2559)
         );
  NOR3_X2 U3516 ( .A1(fract_denorm[80]), .A2(fract_denorm[81]), .A3(
        fract_denorm[79]), .ZN(n2736) );
  OAI21_X2 U3517 ( .B1(n6424), .B2(n6423), .A(n2600), .ZN(n2594) );
  AOI21_X2 U3518 ( .B1(n6336), .B2(n2596), .A(n2597), .ZN(n2595) );
  NAND3_X2 U3519 ( .A1(n6377), .A2(n6379), .A3(n6376), .ZN(n2596) );
  NOR3_X2 U3520 ( .A1(n2598), .A2(n6359), .A3(n2599), .ZN(n2597) );
  AOI211_X2 U3521 ( .C1(fract_denorm[81]), .C2(n6325), .A(n2563), .B(n2573), 
        .ZN(n2572) );
  NAND3_X2 U3522 ( .A1(n6409), .A2(n2711), .A3(n2542), .ZN(n2585) );
  NAND3_X2 U3523 ( .A1(n6416), .A2(n2593), .A3(n2555), .ZN(n2609) );
  NOR3_X2 U3524 ( .A1(fract_denorm[67]), .A2(fract_denorm[68]), .A3(n6396), 
        .ZN(n2646) );
  NOR3_X2 U3525 ( .A1(n2632), .A2(n2696), .A3(n2697), .ZN(n2694) );
  NAND3_X2 U3526 ( .A1(n2707), .A2(fract_denorm[92]), .A3(n6338), .ZN(n2703)
         );
  NOR3_X2 U3527 ( .A1(n2588), .A2(n2625), .A3(n2554), .ZN(n2704) );
  NAND3_X2 U3528 ( .A1(n2708), .A2(n6427), .A3(n2639), .ZN(n2702) );
  NAND3_X2 U3529 ( .A1(n2670), .A2(n6415), .A3(n2555), .ZN(n2607) );
  NOR3_X2 U3530 ( .A1(n6372), .A2(n6370), .A3(n6326), .ZN(n2579) );
  NOR3_X2 U3531 ( .A1(fract_denorm[72]), .A2(fract_denorm[73]), .A3(
        fract_denorm[71]), .ZN(n2661) );
  NOR3_X2 U3532 ( .A1(n6430), .A2(n6431), .A3(n6432), .ZN(n2669) );
  OAI21_X2 U3533 ( .B1(sign), .B2(n3862), .A(n3863), .ZN(n3739) );
  AOI21_X2 U3534 ( .B1(n3880), .B2(n3297), .A(n3881), .ZN(n3862) );
  AOI211_X2 U3535 ( .C1(n3867), .C2(n3868), .A(opas_r2), .B(n4656), .ZN(n3864)
         );
  NAND3_X2 U3536 ( .A1(n3174), .A2(n2752), .A3(n2663), .ZN(n2697) );
  NOR3_X2 U3537 ( .A1(fract_denorm[69]), .A2(fract_denorm[70]), .A3(n6398), 
        .ZN(n2759) );
  NOR3_X2 U3538 ( .A1(fract_denorm[85]), .A2(fract_denorm[86]), .A3(n6378), 
        .ZN(n2760) );
  NOR3_X2 U3539 ( .A1(fract_denorm[56]), .A2(fract_denorm[57]), .A3(
        fract_denorm[55]), .ZN(n2750) );
  NOR3_X2 U3540 ( .A1(fract_denorm[88]), .A2(fract_denorm[89]), .A3(
        fract_denorm[87]), .ZN(n2749) );
  NOR3_X2 U3541 ( .A1(n6423), .A2(n6424), .A3(n6425), .ZN(n2660) );
  NAND3_X2 U3542 ( .A1(n3178), .A2(n2762), .A3(n2695), .ZN(n2635) );
  NOR3_X2 U3543 ( .A1(n2671), .A2(n2771), .A3(n3912), .ZN(n3968) );
  NAND3_X2 U3544 ( .A1(n2644), .A2(n6402), .A3(n6336), .ZN(n2642) );
  NOR3_X2 U3545 ( .A1(n2589), .A2(n6324), .A3(n2557), .ZN(n2727) );
  NAND3_X2 U3546 ( .A1(n6344), .A2(n2724), .A3(n2630), .ZN(n2723) );
  OAI21_X2 U3547 ( .B1(n3865), .B2(n4355), .A(n3866), .ZN(n3853) );
  AOI21_X2 U3548 ( .B1(n3910), .B2(n3911), .A(n3865), .ZN(n3854) );
  NOR3_X2 U3549 ( .A1(remainder[94]), .A2(remainder[96]), .A3(remainder[95]), 
        .ZN(n4165) );
  NOR3_X2 U3550 ( .A1(remainder[88]), .A2(remainder[8]), .A3(remainder[89]), 
        .ZN(n4163) );
  NOR3_X2 U3551 ( .A1(remainder[0]), .A2(remainder[101]), .A3(remainder[100]), 
        .ZN(n4171) );
  NOR3_X2 U3552 ( .A1(remainder[102]), .A2(remainder[104]), .A3(remainder[103]), .ZN(n4172) );
  NOR3_X2 U3553 ( .A1(remainder[105]), .A2(remainder[107]), .A3(remainder[106]), .ZN(n4173) );
  NOR3_X2 U3554 ( .A1(remainder[14]), .A2(remainder[16]), .A3(remainder[15]), 
        .ZN(n4175) );
  NOR3_X2 U3555 ( .A1(remainder[20]), .A2(remainder[22]), .A3(remainder[21]), 
        .ZN(n4177) );
  NOR3_X2 U3556 ( .A1(remainder[27]), .A2(remainder[29]), .A3(remainder[28]), 
        .ZN(n4179) );
  NOR3_X2 U3557 ( .A1(remainder[2]), .A2(remainder[31]), .A3(remainder[30]), 
        .ZN(n4180) );
  NOR3_X2 U3558 ( .A1(remainder[32]), .A2(remainder[34]), .A3(remainder[33]), 
        .ZN(n4181) );
  NOR3_X2 U3559 ( .A1(remainder[39]), .A2(remainder[40]), .A3(remainder[3]), 
        .ZN(n4183) );
  NOR3_X2 U3560 ( .A1(remainder[45]), .A2(remainder[47]), .A3(remainder[46]), 
        .ZN(n4185) );
  NOR3_X2 U3561 ( .A1(remainder[57]), .A2(remainder[59]), .A3(remainder[58]), 
        .ZN(n4153) );
  NOR3_X2 U3562 ( .A1(remainder[63]), .A2(remainder[65]), .A3(remainder[64]), 
        .ZN(n4155) );
  NOR3_X2 U3563 ( .A1(remainder[6]), .A2(remainder[71]), .A3(remainder[70]), 
        .ZN(n4157) );
  NOR3_X2 U3564 ( .A1(remainder[76]), .A2(remainder[78]), .A3(remainder[77]), 
        .ZN(n4159) );
  NOR3_X2 U3565 ( .A1(remainder[79]), .A2(remainder[80]), .A3(remainder[7]), 
        .ZN(n4160) );
  NOR3_X2 U3566 ( .A1(remainder[81]), .A2(remainder[83]), .A3(remainder[82]), 
        .ZN(n4161) );
  NAND3_X2 U3567 ( .A1(n2479), .A2(n4452), .A3(n3487), .ZN(n3486) );
  AOI21_X2 U3568 ( .B1(exp_ovf_r[0]), .B2(n3488), .A(n3489), .ZN(n3487) );
  OAI21_X2 U3569 ( .B1(n2480), .B2(n3494), .A(n3495), .ZN(n3493) );
  NOR3_X2 U3570 ( .A1(n6468), .A2(n4315), .A3(exp_r[1]), .ZN(n3497) );
  OAI21_X2 U3571 ( .B1(n3532), .B2(u4_N6278), .A(n3488), .ZN(n3531) );
  NOR2_X2 U3572 ( .A1(n3488), .A2(n3500), .ZN(n3491) );
  AOI222_X1 U3573 ( .A1(u4_N6284), .A2(u4_N6283), .B1(n3501), .B2(n3502), .C1(
        n3503), .C2(n3495), .ZN(n3500) );
  NAND3_X2 U3574 ( .A1(opb_dn), .A2(n4271), .A3(u4_N6194), .ZN(n3783) );
  AOI21_X2 U3575 ( .B1(n3771), .B2(n3787), .A(n2480), .ZN(n3789) );
  NAND3_X2 U3576 ( .A1(n4353), .A2(n4656), .A3(n4281), .ZN(n3861) );
  OAI21_X2 U3577 ( .B1(n6465), .B2(n4656), .A(n3556), .ZN(n3788) );
  NAND3_X2 U3578 ( .A1(n4403), .A2(n4338), .A3(n4306), .ZN(n3361) );
  NAND3_X2 U3579 ( .A1(n3734), .A2(n3557), .A3(n3735), .ZN(n3733) );
  OAI21_X2 U3580 ( .B1(n3737), .B2(n3477), .A(n3734), .ZN(n3732) );
  NOR3_X2 U3581 ( .A1(n2439), .A2(n6094), .A3(n3736), .ZN(n3735) );
  NOR2_X2 U3582 ( .A1(exp_ovf_r[0]), .A2(exp_ovf_r[1]), .ZN(n3771) );
  OAI21_X2 U3583 ( .B1(exp_ovf_r[1]), .B2(n3551), .A(n3783), .ZN(n3773) );
  NOR3_X2 U3584 ( .A1(n3618), .A2(n3396), .A3(n3398), .ZN(n3746) );
  NAND3_X2 U3585 ( .A1(n3394), .A2(n3395), .A3(n3393), .ZN(n3748) );
  AOI21_X2 U3586 ( .B1(n3834), .B2(rmode_r3[1]), .A(n3835), .ZN(n3795) );
  OAI22_X2 U3587 ( .A1(u4_N6410), .A2(n3847), .B1(n2441), .B2(n2440), .ZN(
        n3805) );
  NOR2_X2 U3588 ( .A1(n3855), .A2(u4_N6203), .ZN(n3798) );
  NOR2_X2 U3589 ( .A1(n6318), .A2(n3855), .ZN(n3799) );
  NOR2_X2 U3590 ( .A1(n3765), .A2(n3477), .ZN(n3761) );
  NAND3_X2 U3591 ( .A1(exp_ovf_r[1]), .A2(n4356), .A3(n4540), .ZN(n3766) );
  INV_X4 U3592 ( .A(n4631), .ZN(n4616) );
  INV_X4 U3593 ( .A(n4632), .ZN(n4631) );
  INV_X4 U3594 ( .A(n4604), .ZN(n4633) );
  NAND3_X2 U3595 ( .A1(n2969), .A2(n6215), .A3(n2970), .ZN(n2963) );
  OAI21_X2 U3596 ( .B1(n2993), .B2(n2994), .A(n2995), .ZN(n2981) );
  OAI21_X2 U3597 ( .B1(n2983), .B2(n2984), .A(n6222), .ZN(n2982) );
  INV_X4 U3598 ( .A(n4633), .ZN(n4627) );
  NOR3_X2 U3599 ( .A1(u6_N12), .A2(u6_N14), .A3(u6_N13), .ZN(n3104) );
  NOR3_X2 U3600 ( .A1(u6_N18), .A2(u6_N1), .A3(u6_N19), .ZN(n3105) );
  NOR3_X2 U3601 ( .A1(u6_N23), .A2(u6_N25), .A3(u6_N24), .ZN(n3106) );
  NOR2_X2 U3602 ( .A1(fracta_mul[34]), .A2(fracta_mul[35]), .ZN(n3283) );
  NOR3_X2 U3603 ( .A1(n3288), .A2(fracta_mul[7]), .A3(n6302), .ZN(n3267) );
  NOR3_X2 U3604 ( .A1(n6297), .A2(fracta_mul[39]), .A3(n6293), .ZN(n3269) );
  NAND3_X2 U3605 ( .A1(n2434), .A2(n2433), .A3(n6317), .ZN(n2508) );
  AOI222_X1 U3606 ( .A1(u4_div_scht1a[6]), .A2(n2484), .B1(u4_f2i_shft_6_), 
        .B2(n6342), .C1(exp_r[6]), .C2(n2483), .ZN(n2491) );
  AOI21_X2 U3607 ( .B1(n2506), .B2(n6316), .A(n6343), .ZN(n2517) );
  NAND3_X2 U3608 ( .A1(n4540), .A2(n2518), .A3(n2515), .ZN(n2516) );
  INV_X4 U3609 ( .A(n2434), .ZN(n6342) );
  NOR2_X2 U3610 ( .A1(n4289), .A2(n4656), .ZN(n3965) );
  AOI211_X2 U3611 ( .C1(n2542), .C2(n6367), .A(n2590), .B(n2591), .ZN(n2574)
         );
  NOR3_X2 U3612 ( .A1(n6391), .A2(n6389), .A3(n6334), .ZN(n2552) );
  NOR3_X2 U3613 ( .A1(n6396), .A2(n6394), .A3(n6335), .ZN(n2549) );
  AOI211_X2 U3614 ( .C1(n2555), .C2(n6412), .A(n2556), .B(n2557), .ZN(n2544)
         );
  OAI21_X2 U3615 ( .B1(n2558), .B2(n6335), .A(n2559), .ZN(n2556) );
  NOR3_X2 U3616 ( .A1(fract_denorm[70]), .A2(fract_denorm[73]), .A3(
        fract_denorm[72]), .ZN(n2558) );
  NOR3_X2 U3617 ( .A1(n6382), .A2(n6381), .A3(n2642), .ZN(n2625) );
  NOR3_X2 U3618 ( .A1(n6385), .A2(n6383), .A3(n2642), .ZN(n2623) );
  NOR3_X2 U3619 ( .A1(n6375), .A2(n6374), .A3(n2671), .ZN(n2620) );
  NAND3_X2 U3620 ( .A1(n2601), .A2(n2602), .A3(n2603), .ZN(n2570) );
  OAI21_X2 U3621 ( .B1(n6384), .B2(n2642), .A(n2643), .ZN(n2573) );
  NAND3_X2 U3622 ( .A1(n2644), .A2(fract_denorm[82]), .A3(n6336), .ZN(n2643)
         );
  NOR3_X2 U3623 ( .A1(n2632), .A2(n2633), .A3(n2634), .ZN(n2631) );
  AOI21_X2 U3624 ( .B1(n6355), .B2(n6356), .A(n2598), .ZN(n2640) );
  OAI21_X2 U3625 ( .B1(n6390), .B2(n6334), .A(n2645), .ZN(n2564) );
  NAND3_X2 U3626 ( .A1(n2646), .A2(fract_denorm[66]), .A3(n2647), .ZN(n2645)
         );
  NAND3_X2 U3627 ( .A1(n2607), .A2(n2666), .A3(n2667), .ZN(n2649) );
  NOR3_X2 U3628 ( .A1(n2586), .A2(n2623), .A3(n2552), .ZN(n2667) );
  NAND3_X2 U3629 ( .A1(n2669), .A2(n6429), .A3(n2639), .ZN(n2666) );
  AOI211_X2 U3630 ( .C1(n2659), .C2(n6349), .A(n2579), .B(n6331), .ZN(n2658)
         );
  NAND3_X2 U3631 ( .A1(n2663), .A2(n6436), .A3(n6327), .ZN(n2655) );
  NAND3_X2 U3632 ( .A1(n2661), .A2(fract_denorm[70]), .A3(n2647), .ZN(n2657)
         );
  NAND3_X2 U3633 ( .A1(n6352), .A2(n6359), .A3(n6338), .ZN(n2671) );
  NOR3_X2 U3634 ( .A1(n2587), .A2(n2624), .A3(n2553), .ZN(n2734) );
  NOR3_X2 U3635 ( .A1(n2584), .A2(n2622), .A3(n2551), .ZN(n2743) );
  NOR2_X2 U3636 ( .A1(n2641), .A2(n2665), .ZN(n2672) );
  NAND3_X2 U3637 ( .A1(n3180), .A2(n2731), .A3(n2709), .ZN(n2561) );
  NOR3_X2 U3638 ( .A1(n6437), .A2(n6438), .A3(n6439), .ZN(n2663) );
  NOR3_X2 U3639 ( .A1(n6350), .A2(n6351), .A3(n2684), .ZN(n2659) );
  NAND3_X2 U3640 ( .A1(n3176), .A2(n2730), .A3(n2708), .ZN(n2604) );
  NAND3_X2 U3641 ( .A1(n6366), .A2(n2770), .A3(n2542), .ZN(n2632) );
  NOR3_X2 U3642 ( .A1(n6380), .A2(fract_denorm[74]), .A3(n2642), .ZN(n2647) );
  NAND3_X2 U3643 ( .A1(n3879), .A2(n2724), .A3(n2630), .ZN(n2710) );
  NOR2_X2 U3644 ( .A1(n3309), .A2(n4482), .ZN(n3565) );
  NOR2_X2 U3645 ( .A1(n6456), .A2(n3304), .ZN(n3568) );
  NAND3_X2 U3646 ( .A1(n3408), .A2(n3409), .A3(n3407), .ZN(n3589) );
  NAND3_X2 U3647 ( .A1(n3600), .A2(n3422), .A3(n3601), .ZN(n3599) );
  AOI211_X2 U3648 ( .C1(n4656), .C2(opas_r2), .A(n2422), .B(n3548), .ZN(n3547)
         );
  NOR2_X2 U3649 ( .A1(n3539), .A2(n3540), .ZN(n3538) );
  OAI21_X2 U3650 ( .B1(exp_ovf_r[0]), .B2(n3483), .A(n3484), .ZN(n3482) );
  NAND3_X2 U3651 ( .A1(n3485), .A2(n4269), .A3(n3486), .ZN(n3484) );
  NAND3_X2 U3652 ( .A1(n4402), .A2(n4342), .A3(n4311), .ZN(n3375) );
  NAND3_X2 U3653 ( .A1(n4401), .A2(n4341), .A3(n4310), .ZN(n3377) );
  NAND3_X2 U3654 ( .A1(n3338), .A2(n3339), .A3(n3337), .ZN(n3438) );
  NOR3_X2 U3655 ( .A1(n3583), .A2(n3584), .A3(n3585), .ZN(n3397) );
  NAND3_X2 U3656 ( .A1(n3430), .A2(n3431), .A3(n3432), .ZN(n3426) );
  NAND3_X2 U3657 ( .A1(n3415), .A2(n3416), .A3(n3417), .ZN(n3411) );
  NAND3_X2 U3658 ( .A1(n6316), .A2(n3467), .A3(n3468), .ZN(n3320) );
  OAI21_X2 U3659 ( .B1(u4_N6410), .B2(n3454), .A(n6454), .ZN(n3467) );
  NAND3_X2 U3660 ( .A1(n3451), .A2(n3452), .A3(n3453), .ZN(n3447) );
  NOR2_X2 U3661 ( .A1(n4356), .A2(n4452), .ZN(n3556) );
  NAND3_X2 U3662 ( .A1(n2434), .A2(n3741), .A3(n3332), .ZN(n3552) );
  AOI222_X1 U3663 ( .A1(u4_exp_out_8_), .A2(n3829), .B1(n3802), .B2(
        u4_exp_next_mi_8_), .C1(u4_exp_out_pl1_8_), .C2(n3805), .ZN(n3846) );
  AOI222_X1 U3664 ( .A1(u4_exp_out_9_), .A2(n3829), .B1(n3802), .B2(
        u4_exp_next_mi_9_), .C1(u4_exp_out_pl1_9_), .C2(n3805), .ZN(n3839) );
  OAI21_X2 U3665 ( .B1(n3762), .B2(n3757), .A(n3758), .ZN(n3585) );
  OAI21_X2 U3666 ( .B1(n3756), .B2(n3757), .A(n3758), .ZN(n3534) );
  NOR2_X2 U3667 ( .A1(n3760), .A2(n3761), .ZN(n3750) );
  INV_X4 U3668 ( .A(n3760), .ZN(n6315) );
  NOR2_X2 U3669 ( .A1(n4262), .A2(fpu_op_r2[1]), .ZN(n4194) );
  INV_X4 U3670 ( .A(n4628), .ZN(n4623) );
  INV_X4 U3671 ( .A(n4619), .ZN(n4607) );
  INV_X4 U3672 ( .A(n4617), .ZN(n4612) );
  INV_X4 U3673 ( .A(n4629), .ZN(n4622) );
  INV_X4 U3674 ( .A(n4618), .ZN(n4610) );
  INV_X4 U3675 ( .A(n4617), .ZN(n4611) );
  AOI21_X2 U3676 ( .B1(n2981), .B2(n2982), .A(n6221), .ZN(n2949) );
  AOI21_X2 U3677 ( .B1(n2951), .B2(n2952), .A(n2953), .ZN(n2950) );
  INV_X4 U3678 ( .A(n4627), .ZN(n4626) );
  INV_X4 U3679 ( .A(u1_fractb_lt_fracta), .ZN(n4635) );
  NOR3_X2 U3680 ( .A1(fracta_mul[40]), .A2(fracta_mul[41]), .A3(n3243), .ZN(
        n3092) );
  NOR3_X2 U3681 ( .A1(fracta_mul[28]), .A2(fracta_mul[29]), .A3(n3217), .ZN(
        n3091) );
  NOR3_X2 U3682 ( .A1(fracta_mul[46]), .A2(fracta_mul[48]), .A3(fracta_mul[47]), .ZN(n3088) );
  NAND3_X2 U3683 ( .A1(n4272), .A2(n4284), .A3(n4276), .ZN(n3087) );
  NOR3_X2 U3684 ( .A1(n6299), .A2(n6296), .A3(n3090), .ZN(n3083) );
  NOR2_X2 U3685 ( .A1(n3219), .A2(n4367), .ZN(n3256) );
  NOR3_X2 U3686 ( .A1(n6299), .A2(fracta_mul[23]), .A3(n3220), .ZN(n3271) );
  NOR3_X2 U3687 ( .A1(n3204), .A2(n6300), .A3(n4318), .ZN(n3290) );
  NOR3_X2 U3688 ( .A1(n4476), .A2(n3225), .A3(n3204), .ZN(n3258) );
  NOR2_X2 U3689 ( .A1(fracta_mul[10]), .A2(fracta_mul[11]), .ZN(n3245) );
  NAND3_X2 U3690 ( .A1(fracta_mul[9]), .A2(n3245), .A3(n6287), .ZN(n3266) );
  NOR2_X2 U3691 ( .A1(n3206), .A2(n4272), .ZN(n3264) );
  NOR3_X2 U3692 ( .A1(n4371), .A2(n3205), .A3(n3204), .ZN(n3268) );
  NAND3_X2 U3693 ( .A1(fracta_mul[6]), .A2(n3267), .A3(n6288), .ZN(n3236) );
  NAND3_X2 U3694 ( .A1(n4326), .A2(n4368), .A3(n3245), .ZN(n3288) );
  NAND3_X2 U3695 ( .A1(n4372), .A2(n4318), .A3(n3246), .ZN(n3225) );
  NOR3_X2 U3696 ( .A1(fracta_mul[12]), .A2(fracta_mul[13]), .A3(n3225), .ZN(
        n3222) );
  NOR3_X2 U3697 ( .A1(n6302), .A2(fracta_mul[9]), .A3(n4326), .ZN(n3223) );
  NAND3_X2 U3698 ( .A1(n4479), .A2(n4370), .A3(n3261), .ZN(n3217) );
  NAND3_X2 U3699 ( .A1(fracta_mul[40]), .A2(n4472), .A3(n3226), .ZN(n3218) );
  NAND3_X2 U3700 ( .A1(fracta_mul[33]), .A2(n3283), .A3(n3260), .ZN(n3259) );
  NOR3_X2 U3701 ( .A1(fracta_mul[4]), .A2(fracta_mul[5]), .A3(n3205), .ZN(
        n3282) );
  NAND3_X2 U3702 ( .A1(fracta_mul[23]), .A2(n3289), .A3(n6284), .ZN(n3229) );
  AOI211_X2 U3703 ( .C1(fracta_mul[26]), .C2(n6281), .A(n6290), .B(n3270), 
        .ZN(n3230) );
  NAND3_X2 U3704 ( .A1(fracta_mul[24]), .A2(n4473), .A3(n6281), .ZN(n3228) );
  NOR3_X2 U3705 ( .A1(fracta_mul[32]), .A2(fracta_mul[33]), .A3(n6298), .ZN(
        n3261) );
  NOR3_X2 U3706 ( .A1(fracta_mul[36]), .A2(fracta_mul[37]), .A3(n3206), .ZN(
        n3260) );
  NOR3_X2 U3707 ( .A1(n4475), .A2(n3217), .A3(n6279), .ZN(n3257) );
  OAI21_X2 U3708 ( .B1(exp_ovf_r[0]), .B2(n2478), .A(n4452), .ZN(n4141) );
  NOR3_X2 U3709 ( .A1(exp_r[6]), .A2(n4353), .A3(n4281), .ZN(n4142) );
  AOI211_X2 U3710 ( .C1(n2562), .C2(fract_denorm[65]), .A(n2563), .B(n2564), 
        .ZN(n2543) );
  NAND2_X2 U3711 ( .A1(n4269), .A2(n4271), .ZN(n3488) );
  NOR3_X2 U3712 ( .A1(n2641), .A2(n2564), .A3(n2573), .ZN(n2627) );
  NOR2_X2 U3713 ( .A1(n3834), .A2(n4351), .ZN(n3848) );
  OAI21_X2 U3714 ( .B1(opb_dn), .B2(n4398), .A(n3170), .ZN(fract_div_105_) );
  NAND3_X2 U3715 ( .A1(n3488), .A2(n2514), .A3(n4455), .ZN(n2479) );
  OAI21_X2 U3716 ( .B1(n2394), .B2(n3528), .A(n3529), .ZN(n3504) );
  AOI222_X1 U3717 ( .A1(u4_div_exp1_10_), .A2(opb_dn), .B1(u4_exp_out1_mi1[10]), .B2(n2397), .C1(u4_div_exp2_10_), .C2(n2398), .ZN(n3528) );
  OAI21_X2 U3718 ( .B1(fract_denorm[102]), .B2(n6363), .A(n6361), .ZN(n2716)
         );
  NAND3_X2 U3719 ( .A1(fract_denorm[99]), .A2(n4653), .A3(n2761), .ZN(n2755)
         );
  NAND3_X2 U3720 ( .A1(n6346), .A2(n2763), .A3(n2700), .ZN(n2754) );
  NAND3_X2 U3721 ( .A1(n6348), .A2(n2751), .A3(n2659), .ZN(n2747) );
  NOR3_X2 U3722 ( .A1(n2580), .A2(n2619), .A3(n2548), .ZN(n2748) );
  NOR3_X2 U3723 ( .A1(n2578), .A2(n2618), .A3(n2547), .ZN(n2766) );
  NOR3_X2 U3724 ( .A1(n2604), .A2(n6441), .A3(n6332), .ZN(n2600) );
  NOR3_X2 U3725 ( .A1(n2592), .A2(fract_denorm[58]), .A3(n6334), .ZN(n2679) );
  NOR2_X2 U3726 ( .A1(n2710), .A2(n6446), .ZN(n2422) );
  NOR2_X2 U3727 ( .A1(n3468), .A2(n4482), .ZN(n3569) );
  NOR2_X2 U3728 ( .A1(qnan_d), .A2(snan_d), .ZN(n3303) );
  NOR3_X2 U3729 ( .A1(n3485), .A2(n3546), .A3(n3547), .ZN(n3542) );
  OAI21_X2 U3730 ( .B1(n3469), .B2(n3470), .A(n3471), .ZN(n3346) );
  NOR2_X2 U3731 ( .A1(n6458), .A2(ind_d), .ZN(n3314) );
  NOR2_X2 U3732 ( .A1(n6458), .A2(inf_d), .ZN(n3457) );
  NOR2_X2 U3733 ( .A1(inf_mul_r), .A2(inf_mul2), .ZN(n3454) );
  NOR2_X2 U3734 ( .A1(n6456), .A2(opb_00), .ZN(n3459) );
  OAI21_X2 U3735 ( .B1(n3764), .B2(n3757), .A(n3758), .ZN(n3584) );
  OAI21_X2 U3736 ( .B1(n3763), .B2(n3757), .A(n3758), .ZN(n3583) );
  AOI21_X2 U3737 ( .B1(n3759), .B2(n6315), .A(n3750), .ZN(n3396) );
  AOI21_X2 U3738 ( .B1(n3755), .B2(n6315), .A(n3750), .ZN(n3540) );
  AOI21_X2 U3739 ( .B1(n3754), .B2(n6315), .A(n3750), .ZN(n3539) );
  AOI21_X2 U3740 ( .B1(n3753), .B2(n6315), .A(n3750), .ZN(n3615) );
  AOI21_X2 U3741 ( .B1(n3752), .B2(n6315), .A(n3750), .ZN(n3389) );
  AOI21_X2 U3742 ( .B1(n3751), .B2(n6315), .A(n3750), .ZN(n3617) );
  AOI21_X2 U3743 ( .B1(n3749), .B2(n6315), .A(n3750), .ZN(n3388) );
  AOI222_X1 U3744 ( .A1(inf_d), .A2(n6339), .B1(opb_00), .B2(n4540), .C1(n4189), .C2(n6316), .ZN(n4188) );
  NOR2_X2 U3745 ( .A1(u4_N6410), .A2(n3454), .ZN(n4189) );
  INV_X4 U3746 ( .A(n4194), .ZN(n6312) );
  NOR2_X2 U3747 ( .A1(fpu_op_r2[1]), .A2(fpu_op_r2[2]), .ZN(n4254) );
  NOR3_X2 U3748 ( .A1(n6275), .A2(n4598), .A3(n6015), .ZN(n2811) );
  NOR3_X2 U3749 ( .A1(n2803), .A2(n6275), .A3(n4597), .ZN(n2810) );
  NOR2_X2 U3750 ( .A1(n6015), .A2(u1_N46), .ZN(n2809) );
  NOR2_X2 U3751 ( .A1(u2_exp_ovf_d_1_), .A2(n6275), .ZN(n2808) );
  NAND2_X2 U3752 ( .A1(n6015), .A2(n6275), .ZN(n2805) );
  NAND3_X2 U3753 ( .A1(u2_N15), .A2(u2_N14), .A3(u2_N6), .ZN(n2781) );
  NAND3_X2 U3754 ( .A1(n4597), .A2(n6032), .A3(u2_N18), .ZN(n2777) );
  NAND3_X2 U3755 ( .A1(u2_N12), .A2(u2_N11), .A3(u2_N13), .ZN(n2780) );
  NOR2_X2 U3756 ( .A1(opb_r[62]), .A2(opa_r[62]), .ZN(n2782) );
  OAI22_X2 U3757 ( .A1(n4599), .A2(n6032), .B1(n4597), .B2(n6017), .ZN(
        u2_exp_tmp4_10_) );
  NOR3_X2 U3758 ( .A1(opa_r1[54]), .A2(opa_r1[56]), .A3(opa_r1[55]), .ZN(n4250) );
  NAND3_X2 U3759 ( .A1(n4484), .A2(n4381), .A3(n4328), .ZN(n4252) );
  INV_X4 U3760 ( .A(n4648), .ZN(n4647) );
  INV_X4 U3761 ( .A(n4648), .ZN(n4646) );
  NOR2_X2 U3762 ( .A1(u1_fracta_eq_fractb), .A2(n3063), .ZN(n3064) );
  AOI211_X2 U3763 ( .C1(n4494), .C2(ind_d), .A(n6458), .B(n3728), .ZN(n3341)
         );
  NOR3_X2 U3764 ( .A1(n4451), .A2(n4456), .A3(n4358), .ZN(n3079) );
  NAND3_X2 U3765 ( .A1(opa_r[61]), .A2(opa_r[62]), .A3(opa_r[60]), .ZN(n3081)
         );
  NOR3_X2 U3766 ( .A1(n4457), .A2(n4359), .A3(n4321), .ZN(n3076) );
  NAND3_X2 U3767 ( .A1(opb_r[61]), .A2(opb_r[62]), .A3(opb_r[60]), .ZN(n3078)
         );
  NOR3_X2 U3768 ( .A1(opa_r[54]), .A2(opa_r[56]), .A3(opa_r[55]), .ZN(n3195)
         );
  NAND3_X2 U3769 ( .A1(n4454), .A2(n4442), .A3(n4453), .ZN(n3197) );
  NOR3_X2 U3770 ( .A1(n3108), .A2(n3109), .A3(n3110), .ZN(n3098) );
  OAI21_X2 U3771 ( .B1(n3279), .B2(n3204), .A(n3266), .ZN(n3278) );
  AOI21_X2 U3772 ( .B1(fracta_mul[17]), .B2(n4369), .A(fracta_mul[19]), .ZN(
        n3279) );
  NOR3_X2 U3773 ( .A1(n4473), .A2(fracta_mul[26]), .A3(n3272), .ZN(n3270) );
  NOR3_X2 U3774 ( .A1(n4472), .A2(n3243), .A3(n6293), .ZN(n3263) );
  NAND3_X2 U3775 ( .A1(fracta_mul[34]), .A2(n4474), .A3(n3260), .ZN(n3254) );
  NAND3_X2 U3776 ( .A1(n4320), .A2(n4283), .A3(n3271), .ZN(n3204) );
  AOI211_X2 U3777 ( .C1(fracta_mul[2]), .C2(n6301), .A(n3274), .B(n3275), .ZN(
        n3273) );
  AOI21_X2 U3778 ( .B1(n4369), .B2(n4319), .A(fracta_mul[19]), .ZN(n3275) );
  NOR2_X2 U3779 ( .A1(fracta_mul[50]), .A2(fracta_mul[49]), .ZN(n3237) );
  AOI21_X2 U3780 ( .B1(n3240), .B2(fracta_mul[47]), .A(n3290), .ZN(n3285) );
  NOR3_X2 U3781 ( .A1(n3287), .A2(n3258), .A3(n3268), .ZN(n3286) );
  NOR3_X2 U3782 ( .A1(fracta_mul[48]), .A2(fracta_mul[51]), .A3(n6296), .ZN(
        n3240) );
  NAND3_X2 U3783 ( .A1(n3207), .A2(n3238), .A3(n3239), .ZN(n3233) );
  NOR3_X2 U3784 ( .A1(fracta_mul[44]), .A2(fracta_mul[45]), .A3(n3219), .ZN(
        n3226) );
  AOI211_X2 U3785 ( .C1(fracta_mul[10]), .C2(n3222), .A(n3223), .B(n3224), 
        .ZN(n3221) );
  NOR3_X2 U3786 ( .A1(n4374), .A2(fracta_mul[13]), .A3(n3225), .ZN(n3224) );
  NAND3_X2 U3787 ( .A1(fracta_mul[3]), .A2(n3282), .A3(n6288), .ZN(n3280) );
  NOR3_X2 U3788 ( .A1(n3204), .A2(fracta_mul[5]), .A3(n3205), .ZN(n3201) );
  NOR2_X2 U3789 ( .A1(n3203), .A2(n6279), .ZN(n3202) );
  NOR3_X2 U3790 ( .A1(fracta_mul[32]), .A2(fracta_mul[34]), .A3(fracta_mul[28]), .ZN(n3203) );
  NOR3_X2 U3791 ( .A1(n3206), .A2(fracta_mul[37]), .A3(n4276), .ZN(n3200) );
  NAND3_X2 U3792 ( .A1(n3228), .A2(n3229), .A3(n3230), .ZN(n3208) );
  NOR3_X2 U3793 ( .A1(n3265), .A2(n3257), .A3(n3291), .ZN(n3198) );
  INV_X4 U3794 ( .A(n3893), .ZN(n4585) );
  NOR2_X2 U3795 ( .A1(u4_N5904), .A2(n3958), .ZN(n3893) );
  NOR3_X2 U3796 ( .A1(n6309), .A2(u4_f2i_shft_9_), .A3(u4_f2i_shft_10_), .ZN(
        n3957) );
  AOI222_X1 U3797 ( .A1(n2483), .A2(n6468), .B1(n2484), .B2(n3960), .C1(n3961), 
        .C2(n2485), .ZN(n3959) );
  INV_X4 U3798 ( .A(n4584), .ZN(n4583) );
  INV_X4 U3799 ( .A(n4585), .ZN(n4584) );
  INV_X4 U3800 ( .A(n4349), .ZN(n4600) );
  NOR2_X2 U3801 ( .A1(n2514), .A2(exp_ovf_r[1]), .ZN(n2480) );
  OAI21_X2 U3802 ( .B1(n4542), .B2(n3522), .A(n3523), .ZN(n2427) );
  AOI222_X1 U3803 ( .A1(u4_div_exp1_8_), .A2(opb_dn), .B1(u4_exp_out1_mi1[8]), 
        .B2(n2397), .C1(u4_div_exp2_8_), .C2(n2398), .ZN(n3522) );
  OAI21_X2 U3804 ( .B1(n4542), .B2(n3526), .A(n3527), .ZN(n2423) );
  AOI222_X1 U3805 ( .A1(u4_div_exp1_7_), .A2(opb_dn), .B1(u4_exp_out1_mi1[7]), 
        .B2(n2397), .C1(u4_div_exp2_7_), .C2(n2398), .ZN(n3526) );
  OAI21_X2 U3806 ( .B1(n2394), .B2(n3515), .A(n3516), .ZN(n2413) );
  AOI222_X1 U3807 ( .A1(u4_div_exp1_3_), .A2(opb_dn), .B1(u4_exp_out1_mi1[3]), 
        .B2(n2397), .C1(u4_div_exp2_3_), .C2(n2398), .ZN(n3515) );
  OAI21_X2 U3808 ( .B1(n2394), .B2(n3519), .A(n3520), .ZN(n2410) );
  AOI222_X1 U3809 ( .A1(u4_div_exp1_2_), .A2(opb_dn), .B1(u4_exp_out1_mi1[2]), 
        .B2(n2397), .C1(u4_div_exp2_2_), .C2(n2398), .ZN(n3519) );
  NAND3_X2 U3810 ( .A1(fpu_op_r3[0]), .A2(n4400), .A3(n4661), .ZN(n2434) );
  OAI21_X2 U3811 ( .B1(fract_denorm[105]), .B2(n6096), .A(n3964), .ZN(n2438)
         );
  NOR2_X2 U3812 ( .A1(n4452), .A2(n2507), .ZN(n2441) );
  NAND3_X2 U3813 ( .A1(n4274), .A2(n4400), .A3(n4661), .ZN(n2433) );
  INV_X4 U3814 ( .A(n4440), .ZN(n4656) );
  NOR2_X2 U3815 ( .A1(n4355), .A2(n3913), .ZN(n2449) );
  NOR2_X2 U3816 ( .A1(n4540), .A2(n2480), .ZN(n2447) );
  NOR3_X2 U3817 ( .A1(n4355), .A2(n6448), .A3(n2479), .ZN(n2448) );
  OAI21_X2 U3818 ( .B1(n2394), .B2(n3524), .A(n3525), .ZN(n2430) );
  AOI222_X1 U3819 ( .A1(u4_div_exp1_9_), .A2(opb_dn), .B1(u4_exp_out1_mi1[9]), 
        .B2(n2397), .C1(u4_div_exp2_9_), .C2(n2398), .ZN(n3524) );
  OAI21_X2 U3820 ( .B1(n4542), .B2(n3517), .A(n3518), .ZN(n2406) );
  AOI222_X1 U3821 ( .A1(u4_div_exp1_1_), .A2(opb_dn), .B1(u4_exp_out1_mi1[1]), 
        .B2(n2397), .C1(u4_div_exp2_1_), .C2(n2398), .ZN(n3517) );
  OAI21_X2 U3822 ( .B1(n4542), .B2(n2395), .A(n2396), .ZN(n2393) );
  AOI222_X1 U3823 ( .A1(u4_div_exp1_0_), .A2(opb_dn), .B1(u4_exp_out1_mi1[0]), 
        .B2(n2397), .C1(u4_div_exp2_0_), .C2(n2398), .ZN(n2395) );
  NOR2_X2 U3824 ( .A1(n2422), .A2(n2433), .ZN(n2390) );
  OAI21_X2 U3825 ( .B1(n3302), .B2(n3558), .A(n3559), .ZN(N875) );
  OAI21_X2 U3826 ( .B1(n3301), .B2(n3302), .A(n3303), .ZN(n3300) );
  OAI21_X2 U3827 ( .B1(opb_00), .B2(n3304), .A(n4327), .ZN(n3307) );
  NAND3_X2 U3828 ( .A1(n4595), .A2(n3463), .A3(n3457), .ZN(n3462) );
  AOI21_X2 U3829 ( .B1(n3465), .B2(n3466), .A(opa_00), .ZN(n3464) );
  OAI21_X2 U3830 ( .B1(n3386), .B2(n3319), .A(n3387), .ZN(n3345) );
  NAND3_X2 U3831 ( .A1(n3314), .A2(n4595), .A3(inf_d), .ZN(n3313) );
  AOI21_X2 U3832 ( .B1(n3316), .B2(n4291), .A(n3317), .ZN(n3312) );
  NOR2_X2 U3833 ( .A1(n6310), .A2(n3330), .ZN(N794) );
  NOR2_X2 U3834 ( .A1(n6310), .A2(n3329), .ZN(N795) );
  NOR2_X2 U3835 ( .A1(n4545), .A2(n3437), .ZN(N796) );
  NOR2_X2 U3836 ( .A1(n6310), .A2(n3582), .ZN(N797) );
  NOR2_X2 U3837 ( .A1(n4545), .A2(n3581), .ZN(N798) );
  NOR2_X2 U3838 ( .A1(n4545), .A2(n3340), .ZN(N799) );
  NOR2_X2 U3839 ( .A1(n4545), .A2(n3339), .ZN(N800) );
  NOR2_X2 U3840 ( .A1(n4545), .A2(n3338), .ZN(N801) );
  NOR2_X2 U3841 ( .A1(n4545), .A2(n3337), .ZN(N802) );
  NOR2_X2 U3842 ( .A1(n4545), .A2(n3580), .ZN(N803) );
  NOR2_X2 U3843 ( .A1(n4545), .A2(n3579), .ZN(N804) );
  NOR2_X2 U3844 ( .A1(n4545), .A2(n3578), .ZN(N805) );
  NOR2_X2 U3845 ( .A1(n4545), .A2(n3446), .ZN(N806) );
  NOR2_X2 U3846 ( .A1(n4545), .A2(n3445), .ZN(N807) );
  NOR2_X2 U3847 ( .A1(n4545), .A2(n3444), .ZN(N808) );
  NOR2_X2 U3848 ( .A1(n4544), .A2(n3443), .ZN(N809) );
  NOR2_X2 U3849 ( .A1(n4544), .A2(n3595), .ZN(N810) );
  NOR2_X2 U3850 ( .A1(n4544), .A2(n3594), .ZN(N811) );
  NOR2_X2 U3851 ( .A1(n4544), .A2(n3593), .ZN(N812) );
  NOR2_X2 U3852 ( .A1(n4544), .A2(n3452), .ZN(N813) );
  NOR2_X2 U3853 ( .A1(n4544), .A2(n3451), .ZN(N814) );
  NOR2_X2 U3854 ( .A1(n4544), .A2(n3453), .ZN(N815) );
  NOR2_X2 U3855 ( .A1(n4544), .A2(n3592), .ZN(N816) );
  NOR2_X2 U3856 ( .A1(n4544), .A2(n3591), .ZN(N817) );
  NOR2_X2 U3857 ( .A1(n4544), .A2(n3590), .ZN(N818) );
  NOR2_X2 U3858 ( .A1(n4544), .A2(n3410), .ZN(N819) );
  NOR2_X2 U3859 ( .A1(n4544), .A2(n3409), .ZN(N820) );
  NOR2_X2 U3860 ( .A1(n4543), .A2(n3408), .ZN(N821) );
  NOR2_X2 U3861 ( .A1(n4545), .A2(n3407), .ZN(N822) );
  NOR2_X2 U3862 ( .A1(n4545), .A2(n3607), .ZN(N823) );
  NOR2_X2 U3863 ( .A1(n4543), .A2(n3606), .ZN(N824) );
  NOR2_X2 U3864 ( .A1(n4543), .A2(n3605), .ZN(N825) );
  NOR2_X2 U3865 ( .A1(n4545), .A2(n3416), .ZN(N826) );
  NOR2_X2 U3866 ( .A1(n4544), .A2(n3415), .ZN(N827) );
  NOR2_X2 U3867 ( .A1(n4543), .A2(n3417), .ZN(N828) );
  NOR2_X2 U3868 ( .A1(n4544), .A2(n3604), .ZN(N829) );
  NOR2_X2 U3869 ( .A1(n4544), .A2(n3603), .ZN(N830) );
  NOR2_X2 U3870 ( .A1(n4545), .A2(n3602), .ZN(N831) );
  NOR2_X2 U3871 ( .A1(n4543), .A2(n3425), .ZN(N832) );
  NOR2_X2 U3872 ( .A1(n4543), .A2(n3424), .ZN(N833) );
  NOR2_X2 U3873 ( .A1(n4544), .A2(n3423), .ZN(N834) );
  NOR2_X2 U3874 ( .A1(n4543), .A2(n3422), .ZN(N835) );
  NOR2_X2 U3875 ( .A1(n4543), .A2(n3600), .ZN(N836) );
  NOR2_X2 U3876 ( .A1(n4543), .A2(n3601), .ZN(N837) );
  NOR2_X2 U3877 ( .A1(n4543), .A2(n3614), .ZN(N838) );
  NOR2_X2 U3878 ( .A1(n4543), .A2(n3431), .ZN(N839) );
  NOR2_X2 U3879 ( .A1(n4543), .A2(n3430), .ZN(N840) );
  NOR2_X2 U3880 ( .A1(n4543), .A2(n3432), .ZN(N841) );
  NOR2_X2 U3881 ( .A1(n4543), .A2(n3613), .ZN(N842) );
  NOR2_X2 U3882 ( .A1(n4543), .A2(n3612), .ZN(N843) );
  NOR2_X2 U3883 ( .A1(n4543), .A2(n3611), .ZN(N844) );
  AOI21_X2 U3884 ( .B1(n3457), .B2(n3458), .A(n3459), .ZN(n3455) );
  NOR3_X2 U3885 ( .A1(opb_r[54]), .A2(opb_r[56]), .A3(opb_r[55]), .ZN(n3093)
         );
  NAND3_X2 U3886 ( .A1(n4399), .A2(n4340), .A3(n4296), .ZN(n3095) );
  NAND3_X2 U3887 ( .A1(exp_mul[6]), .A2(exp_mul[5]), .A3(exp_mul[7]), .ZN(
        n3294) );
  NOR3_X2 U3888 ( .A1(n4487), .A2(n4383), .A3(n4330), .ZN(n3295) );
  NAND3_X2 U3889 ( .A1(n6016), .A2(n4597), .A3(n2782), .ZN(n2832) );
  AOI21_X2 U3890 ( .B1(n2801), .B2(n2802), .A(n4458), .ZN(u2_exp_ovf_d_0_) );
  NOR2_X2 U3891 ( .A1(n2772), .A2(n6274), .ZN(u2_underflow_d[2]) );
  OAI21_X2 U3892 ( .B1(n4597), .B2(n2833), .A(n2834), .ZN(u2_N114) );
  OAI21_X2 U3893 ( .B1(n4191), .B2(n4380), .A(n4203), .ZN(N710) );
  OAI21_X2 U3894 ( .B1(n4191), .B2(n4488), .A(n4202), .ZN(N711) );
  NOR2_X2 U3895 ( .A1(n3059), .A2(n6262), .ZN(u1_N62) );
  NOR2_X2 U3896 ( .A1(n3059), .A2(n3050), .ZN(u1_N61) );
  NOR2_X2 U3897 ( .A1(n3059), .A2(n3051), .ZN(u1_N60) );
  NOR2_X2 U3898 ( .A1(n3059), .A2(n6265), .ZN(u1_N59) );
  NOR2_X2 U3899 ( .A1(n3059), .A2(n6266), .ZN(u1_N58) );
  NOR2_X2 U3900 ( .A1(n3059), .A2(n6267), .ZN(u1_N57) );
  NOR2_X2 U3901 ( .A1(n3059), .A2(n6268), .ZN(u1_N56) );
  NOR2_X2 U3902 ( .A1(n3059), .A2(n6269), .ZN(u1_N55) );
  NOR2_X2 U3903 ( .A1(n3059), .A2(n6270), .ZN(u1_N54) );
  NOR2_X2 U3904 ( .A1(n3059), .A2(n6271), .ZN(u1_N53) );
  NOR2_X2 U3905 ( .A1(n3059), .A2(n6272), .ZN(u1_N52) );
  OAI21_X2 U3906 ( .B1(n3060), .B2(n4495), .A(n3061), .ZN(u1_N229) );
  OAI21_X2 U3907 ( .B1(n3062), .B2(n4492), .A(u1_signa_r), .ZN(n3061) );
  NOR3_X2 U3908 ( .A1(n3063), .A2(u1_fracta_lt_fractb), .A3(
        u1_fracta_eq_fractb), .ZN(n3062) );
  NOR2_X2 U3909 ( .A1(n4661), .A2(n3341), .ZN(N904) );
  NOR2_X2 U3910 ( .A1(n3071), .A2(n3070), .ZN(u0_N6) );
  NOR2_X2 U3911 ( .A1(fracta_mul[51]), .A2(n3073), .ZN(u0_N4) );
  NOR3_X2 U3912 ( .A1(n4493), .A2(opa_nan), .A3(n3296), .ZN(N912) );
  NOR2_X2 U3913 ( .A1(n4267), .A2(n3075), .ZN(u0_N10) );
  NOR2_X2 U3914 ( .A1(n4268), .A2(n3074), .ZN(u0_N11) );
  NOR2_X2 U3915 ( .A1(n3072), .A2(u6_N51), .ZN(n4268) );
  AOI21_X2 U3916 ( .B1(fracta_mul[49]), .B2(n4480), .A(n3209), .ZN(n3276) );
  NOR2_X2 U3917 ( .A1(n3273), .A2(n3204), .ZN(n3249) );
  AOI211_X2 U3918 ( .C1(n3240), .C2(fracta_mul[46]), .A(n3241), .B(n3242), 
        .ZN(n3231) );
  AOI211_X2 U3919 ( .C1(n3226), .C2(fracta_mul[42]), .A(n3227), .B(n3208), 
        .ZN(n3212) );
  NOR3_X2 U3920 ( .A1(n3219), .A2(fracta_mul[45]), .A3(n4277), .ZN(n3215) );
  INV_X4 U3921 ( .A(n4583), .ZN(n4579) );
  INV_X4 U3922 ( .A(n4585), .ZN(n4580) );
  INV_X4 U3923 ( .A(n4583), .ZN(n4581) );
  INV_X4 U3924 ( .A(n4585), .ZN(n4582) );
  INV_X4 U3925 ( .A(n4583), .ZN(n4578) );
  NAND2_X2 U3926 ( .A1(n2480), .A2(n4355), .ZN(n2442) );
  OAI21_X2 U3927 ( .B1(n4542), .B2(n3513), .A(n3514), .ZN(n3512) );
  AOI222_X1 U3928 ( .A1(u4_div_exp1_6_), .A2(opb_dn), .B1(u4_exp_out1_mi1[6]), 
        .B2(n2397), .C1(u4_div_exp2_6_), .C2(n2398), .ZN(n3513) );
  OAI21_X2 U3929 ( .B1(n2394), .B2(n3507), .A(n3508), .ZN(n3506) );
  AOI222_X1 U3930 ( .A1(u4_div_exp1_5_), .A2(opb_dn), .B1(u4_exp_out1_mi1[5]), 
        .B2(n2397), .C1(u4_div_exp2_5_), .C2(n2398), .ZN(n3507) );
  OAI21_X2 U3931 ( .B1(n2394), .B2(n3510), .A(n3511), .ZN(n3509) );
  AOI222_X1 U3932 ( .A1(u4_div_exp1_4_), .A2(opb_dn), .B1(u4_exp_out1_mi1[4]), 
        .B2(n2397), .C1(u4_div_exp2_4_), .C2(n2398), .ZN(n3510) );
  INV_X4 U3933 ( .A(n2401), .ZN(n2408) );
  NOR3_X2 U3934 ( .A1(n2434), .A2(n6309), .A3(n2435), .ZN(n2400) );
  NAND3_X2 U3935 ( .A1(n2436), .A2(n2433), .A3(n2437), .ZN(n2399) );
  AOI21_X2 U3936 ( .B1(n6316), .B2(n2438), .A(n2439), .ZN(n2437) );
  NAND3_X2 U3937 ( .A1(n2440), .A2(n4356), .A3(n2441), .ZN(n2436) );
  AOI222_X1 U3938 ( .A1(u4_fi_ldz_2a_0_), .A2(n2390), .B1(n2391), .B2(n6094), 
        .C1(n4540), .C2(n2393), .ZN(n2389) );
  NOR3_X2 U3939 ( .A1(u4_N5945), .A2(u4_N5947), .A3(u4_N5946), .ZN(n3932) );
  NOR3_X2 U3940 ( .A1(u4_N5952), .A2(u4_N5954), .A3(u4_N5953), .ZN(n3934) );
  NOR3_X2 U3941 ( .A1(u4_N5932), .A2(u4_N5934), .A3(u4_N5933), .ZN(n3928) );
  NOR3_X2 U3942 ( .A1(u4_N5935), .A2(u4_N5937), .A3(u4_N5936), .ZN(n3929) );
  NOR3_X2 U3943 ( .A1(u4_N5938), .A2(u4_N5940), .A3(u4_N5939), .ZN(n3930) );
  NOR3_X2 U3944 ( .A1(u4_N5919), .A2(u4_N5921), .A3(u4_N5920), .ZN(n3924) );
  NOR3_X2 U3945 ( .A1(u4_N5922), .A2(u4_N5924), .A3(u4_N5923), .ZN(n3925) );
  NOR3_X2 U3946 ( .A1(u4_N5925), .A2(u4_N5927), .A3(u4_N5926), .ZN(n3926) );
  NOR3_X2 U3947 ( .A1(u4_N5906), .A2(u4_N5908), .A3(u4_N5907), .ZN(n3920) );
  NOR3_X2 U3948 ( .A1(u4_N5909), .A2(u4_N5911), .A3(u4_N5910), .ZN(n3921) );
  NOR3_X2 U3949 ( .A1(u4_N5912), .A2(u4_N5914), .A3(u4_N5913), .ZN(n3922) );
  INV_X4 U3950 ( .A(n4620), .ZN(n4606) );
  INV_X4 U3951 ( .A(n4650), .ZN(n4642) );
  INV_X4 U3952 ( .A(n4630), .ZN(n4619) );
  INV_X4 U3953 ( .A(n4616), .ZN(n4615) );
  INV_X4 U3954 ( .A(n4569), .ZN(n4566) );
  INV_X4 U3955 ( .A(n4568), .ZN(n4567) );
  INV_X4 U3956 ( .A(n4632), .ZN(n4630) );
  INV_X4 U3957 ( .A(n4660), .ZN(n4659) );
  INV_X4 U3958 ( .A(n4632), .ZN(n4629) );
  AND2_X4 U3959 ( .A1(n3734), .A2(n3742), .ZN(n4278) );
  AND2_X4 U3960 ( .A1(n3734), .A2(n3738), .ZN(n4279) );
  OR2_X4 U3961 ( .A1(n4269), .A2(n3458), .ZN(n4280) );
  INV_X4 U3962 ( .A(n4634), .ZN(n4650) );
  INV_X4 U3963 ( .A(n4635), .ZN(n4634) );
  INV_X4 U3964 ( .A(n4633), .ZN(n4628) );
  INV_X4 U3965 ( .A(n4629), .ZN(n4621) );
  NAND2_X2 U3966 ( .A1(n3732), .A2(n3733), .ZN(n4288) );
  INV_X4 U3967 ( .A(n4565), .ZN(n4564) );
  INV_X4 U3968 ( .A(n4634), .ZN(n4645) );
  INV_X4 U3969 ( .A(n4634), .ZN(n4644) );
  INV_X4 U3970 ( .A(n4634), .ZN(n4643) );
  NOR2_X2 U3971 ( .A1(n4271), .A2(n4269), .ZN(n2394) );
  INV_X4 U3972 ( .A(n4541), .ZN(n4542) );
  INV_X4 U3973 ( .A(n4631), .ZN(n4618) );
  NAND2_X2 U3974 ( .A1(n4187), .A2(n2433), .ZN(n3619) );
  AND2_X4 U3975 ( .A1(n6312), .A2(n6313), .ZN(n4293) );
  INV_X4 U3976 ( .A(n4291), .ZN(n4661) );
  NOR3_X2 U3977 ( .A1(u4_N6172), .A2(u4_N6171), .A3(n4271), .ZN(n2398) );
  INV_X4 U3978 ( .A(n4280), .ZN(n4572) );
  INV_X4 U3979 ( .A(n3973), .ZN(n4569) );
  INV_X4 U3980 ( .A(n4650), .ZN(n4639) );
  INV_X4 U3981 ( .A(n4644), .ZN(n4637) );
  INV_X4 U3982 ( .A(n4645), .ZN(n4636) );
  AND3_X4 U3983 ( .A1(n4194), .A2(n6313), .A3(N396), .ZN(n4302) );
  OR2_X4 U3984 ( .A1(n6312), .A2(n6313), .ZN(n4304) );
  NOR2_X2 U3985 ( .A1(n3458), .A2(opb_dn), .ZN(n4309) );
  INV_X4 U3986 ( .A(n4280), .ZN(n4570) );
  INV_X4 U3987 ( .A(n3956), .ZN(n4576) );
  NOR2_X2 U3988 ( .A1(n3488), .A2(n2480), .ZN(n2397) );
  INV_X4 U3989 ( .A(n4650), .ZN(n4641) );
  INV_X4 U3990 ( .A(n4650), .ZN(n4640) );
  INV_X4 U3991 ( .A(n4650), .ZN(n4638) );
  INV_X4 U3992 ( .A(u2_N157), .ZN(n4601) );
  INV_X8 U3993 ( .A(n4603), .ZN(n4602) );
  INV_X4 U3994 ( .A(u2_N157), .ZN(n4603) );
  INV_X4 U3995 ( .A(n4631), .ZN(n4617) );
  INV_X4 U3996 ( .A(n4302), .ZN(n4556) );
  INV_X4 U3997 ( .A(n4302), .ZN(n4554) );
  INV_X4 U3998 ( .A(n4302), .ZN(n4555) );
  INV_X4 U3999 ( .A(n3619), .ZN(n4545) );
  INV_X4 U4000 ( .A(n3619), .ZN(n4543) );
  INV_X4 U4001 ( .A(n3619), .ZN(n4544) );
  INV_X4 U4002 ( .A(n4379), .ZN(n4598) );
  INV_X4 U4003 ( .A(n4598), .ZN(n4597) );
  INV_X4 U4004 ( .A(n4562), .ZN(n4561) );
  NOR2_X2 U4005 ( .A1(n6312), .A2(n4190), .ZN(n4197) );
  OR2_X4 U4006 ( .A1(n4720), .A2(u4_exp_out_4_), .ZN(n4337) );
  OR2_X4 U4007 ( .A1(n4713), .A2(u4_sub_468_A_4_), .ZN(n4339) );
  NOR2_X2 U4008 ( .A1(fpu_op_r3[1]), .A2(n4661), .ZN(n3315) );
  INV_X4 U4009 ( .A(n4278), .ZN(n4593) );
  INV_X4 U4010 ( .A(n4288), .ZN(n4586) );
  INV_X4 U4011 ( .A(n4280), .ZN(n4574) );
  INV_X4 U4012 ( .A(n4280), .ZN(n4573) );
  INV_X4 U4013 ( .A(n4309), .ZN(n4565) );
  INV_X4 U4014 ( .A(n4291), .ZN(n4662) );
  INV_X4 U4015 ( .A(n4653), .ZN(n4652) );
  INV_X4 U4016 ( .A(n4652), .ZN(n4654) );
  INV_X4 U4017 ( .A(fract_denorm[105]), .ZN(n4653) );
  INV_X4 U4018 ( .A(n3973), .ZN(n4568) );
  OR2_X4 U4019 ( .A1(n4692), .A2(exp_r[6]), .ZN(n4354) );
  INV_X4 U4020 ( .A(n4316), .ZN(n4655) );
  OR2_X4 U4021 ( .A1(n3458), .A2(n4661), .ZN(n4355) );
  INV_X4 U4022 ( .A(n4651), .ZN(n4648) );
  INV_X4 U4023 ( .A(n4634), .ZN(n4651) );
  NAND4_X2 U4024 ( .A1(n2712), .A2(n2713), .A3(n2714), .A4(n2715), .ZN(
        u4_fi_ldz_2a_0_) );
  OR2_X4 U4025 ( .A1(n4679), .A2(u2_exp_tmp4_4_), .ZN(n4378) );
  NAND3_X2 U4026 ( .A1(fpu_op_r1[0]), .A2(n4377), .A3(fpu_op_r1[1]), .ZN(n4379) );
  INV_X4 U4027 ( .A(n4191), .ZN(n4562) );
  INV_X4 U4028 ( .A(n4304), .ZN(n4552) );
  INV_X4 U4029 ( .A(n4293), .ZN(n4558) );
  INV_X4 U4030 ( .A(n4293), .ZN(n4557) );
  INV_X4 U4031 ( .A(n4305), .ZN(n4657) );
  INV_X4 U4032 ( .A(n4305), .ZN(n4658) );
  NOR2_X2 U4033 ( .A1(n2518), .A2(n4355), .ZN(n2483) );
  INV_X4 U4034 ( .A(n4279), .ZN(n4590) );
  INV_X4 U4035 ( .A(n4279), .ZN(n4591) );
  INV_X4 U4036 ( .A(n4279), .ZN(n4589) );
  INV_X4 U4037 ( .A(n4278), .ZN(n4592) );
  INV_X4 U4038 ( .A(n4278), .ZN(n4594) );
  INV_X4 U4039 ( .A(n4288), .ZN(n4587) );
  INV_X4 U4040 ( .A(n4288), .ZN(n4588) );
  INV_X4 U4041 ( .A(n3315), .ZN(n4596) );
  INV_X4 U4042 ( .A(n4596), .ZN(n4595) );
  NAND4_X2 U4043 ( .A1(n2626), .A2(n2627), .A3(n2628), .A4(n2629), .ZN(
        u4_fi_ldz_3_) );
  INV_X4 U4044 ( .A(n4280), .ZN(n4571) );
  INV_X4 U4045 ( .A(n4280), .ZN(n4575) );
  INV_X4 U4046 ( .A(n4565), .ZN(n4563) );
  NAND4_X2 U4047 ( .A1(n2565), .A2(n2566), .A3(n2567), .A4(n2568), .ZN(
        u4_fi_ldz_4_) );
  NAND4_X2 U4048 ( .A1(n2543), .A2(n2544), .A3(n2545), .A4(n2546), .ZN(
        u4_fi_ldz_5_) );
  INV_X4 U4049 ( .A(n3956), .ZN(n4577) );
  NOR2_X2 U4050 ( .A1(n4352), .A2(u4_sub_409_carry[10]), .ZN(n4455) );
  INV_X4 U4051 ( .A(n2394), .ZN(n4541) );
  INV_X4 U4052 ( .A(n4650), .ZN(n4649) );
  INV_X4 U4053 ( .A(n4355), .ZN(n4540) );
  INV_X4 U4054 ( .A(n4630), .ZN(n4620) );
  NAND2_X2 U4055 ( .A1(n4351), .A2(n4441), .ZN(u4_N6410) );
  INV_X4 U4056 ( .A(n2800), .ZN(u2_lt_135_A_0_) );
  INV_X4 U4057 ( .A(n4304), .ZN(n4553) );
  INV_X4 U4058 ( .A(n4304), .ZN(n4550) );
  INV_X4 U4059 ( .A(n4304), .ZN(n4551) );
  INV_X4 U4060 ( .A(n4197), .ZN(n4549) );
  INV_X4 U4061 ( .A(n4549), .ZN(n4546) );
  INV_X4 U4062 ( .A(n4549), .ZN(n4547) );
  INV_X4 U4063 ( .A(n4549), .ZN(n4548) );
  INV_X4 U4064 ( .A(n4293), .ZN(n4559) );
  INV_X4 U4065 ( .A(n4293), .ZN(n4560) );
  INV_X4 U4066 ( .A(n4305), .ZN(n4660) );
  INV_X4 U4067 ( .A(n4379), .ZN(n4599) );
  OAI22_X2 U4068 ( .A1(u4_fi_ldz_2a_6_), .A2(n4812), .B1(u4_fi_ldz_2a_6_), 
        .B2(u4_fi_ldz_2a_5_), .ZN(u4_N6249) );
  OR2_X4 U4069 ( .A1(n4303), .A2(fpu_op_r2[2]), .ZN(n3296) );
  AND2_X4 U4070 ( .A1(n3848), .A2(n2441), .ZN(n3804) );
  AND3_X4 U4071 ( .A1(n6305), .A2(n4355), .A3(n3849), .ZN(n3802) );
  AND3_X4 U4072 ( .A1(u1_N220), .A2(n6099), .A3(u1_N49), .ZN(n3059) );
  AND3_X4 U4073 ( .A1(n6404), .A2(n6403), .A3(n2637), .ZN(n2542) );
  OR4_X4 U4074 ( .A1(n2651), .A2(n2652), .A3(n2653), .A4(n2654), .ZN(
        u4_fi_ldz_2_) );
  AND2_X4 U4075 ( .A1(n2478), .A2(n4540), .ZN(n2446) );
  XNOR2_X1 U4076 ( .A(u4_fi_ldz_6_), .B(u4_sub_463_carry_6_), .ZN(
        u4_fi_ldz_mi22[6]) );
  AND2_X1 U4077 ( .A1(u4_sub_463_carry_5_), .A2(u4_fi_ldz_5_), .ZN(
        u4_sub_463_carry_6_) );
  XOR2_X1 U4078 ( .A(u4_fi_ldz_5_), .B(u4_sub_463_carry_5_), .Z(
        u4_fi_ldz_mi22[5]) );
  AND2_X1 U4079 ( .A1(u4_sub_463_carry_4_), .A2(u4_fi_ldz_4_), .ZN(
        u4_sub_463_carry_5_) );
  XOR2_X1 U4080 ( .A(u4_fi_ldz_4_), .B(u4_sub_463_carry_4_), .Z(
        u4_fi_ldz_mi22[4]) );
  OR2_X1 U4081 ( .A1(u4_fi_ldz_3_), .A2(u4_sub_463_carry_3_), .ZN(
        u4_sub_463_carry_4_) );
  XNOR2_X1 U4082 ( .A(u4_sub_463_carry_3_), .B(u4_fi_ldz_3_), .ZN(
        u4_fi_ldz_mi22[3]) );
  OR2_X1 U4083 ( .A1(u4_fi_ldz_2_), .A2(u4_sub_463_carry_2_), .ZN(
        u4_sub_463_carry_3_) );
  XNOR2_X1 U4084 ( .A(u4_sub_463_carry_2_), .B(u4_fi_ldz_2_), .ZN(
        u4_fi_ldz_mi22[2]) );
  AND2_X1 U4085 ( .A1(u4_fi_ldz_2a_0_), .A2(u4_fi_ldz_1_), .ZN(
        u4_sub_463_carry_2_) );
  XOR2_X1 U4086 ( .A(u4_fi_ldz_1_), .B(u4_fi_ldz_2a_0_), .Z(u4_fi_ldz_mi22[1])
         );
  XOR2_X1 U4087 ( .A(n4656), .B(u4_add_410_carry[10]), .Z(u4_div_shft2[10]) );
  AND2_X1 U4088 ( .A1(n4289), .A2(u4_add_410_carry[9]), .ZN(
        u4_add_410_carry[10]) );
  XOR2_X1 U4089 ( .A(n4289), .B(u4_add_410_carry[9]), .Z(u4_div_shft2[9]) );
  XOR2_X1 U4090 ( .A(n4656), .B(u4_add_411_carry[10]), .Z(u4_div_shft3_10_) );
  AND2_X1 U4091 ( .A1(n4289), .A2(u4_add_411_carry[9]), .ZN(
        u4_add_411_carry[10]) );
  XOR2_X1 U4092 ( .A(n4289), .B(u4_add_411_carry[9]), .Z(u4_div_shft3_9_) );
  XOR2_X1 U4093 ( .A(n4440), .B(u4_sub_412_carry[10]), .Z(u4_div_shft4[10]) );
  AND2_X1 U4094 ( .A1(u4_sub_412_carry[9]), .A2(n4350), .ZN(
        u4_sub_412_carry[10]) );
  XOR2_X1 U4095 ( .A(n4350), .B(u4_sub_412_carry[9]), .Z(u4_div_shft4[9]) );
  XNOR2_X1 U4096 ( .A(n4656), .B(sub_1_root_sub_0_root_u4_add_497_carry[10]), 
        .ZN(u4_ldz_dif_10_) );
  OR2_X1 U4097 ( .A1(n4289), .A2(sub_1_root_sub_0_root_u4_add_497_carry[9]), 
        .ZN(sub_1_root_sub_0_root_u4_add_497_carry[10]) );
  XNOR2_X1 U4098 ( .A(sub_1_root_sub_0_root_u4_add_497_carry[9]), .B(n4289), 
        .ZN(u4_ldz_dif_9_) );
  AND2_X1 U4099 ( .A1(n4353), .A2(u4_add_410_carry[8]), .ZN(
        u4_add_410_carry[9]) );
  XOR2_X1 U4100 ( .A(n4353), .B(u4_add_410_carry[8]), .Z(u4_div_shft2[8]) );
  AND2_X1 U4101 ( .A1(n4353), .A2(u4_add_411_carry[8]), .ZN(
        u4_add_411_carry[9]) );
  XOR2_X1 U4102 ( .A(n4353), .B(u4_add_411_carry[8]), .Z(u4_div_shft3_8_) );
  AND2_X1 U4103 ( .A1(u4_sub_412_carry[8]), .A2(n4439), .ZN(
        u4_sub_412_carry[9]) );
  XOR2_X1 U4104 ( .A(n4439), .B(u4_sub_412_carry[8]), .Z(u4_div_shft4[8]) );
  OR2_X1 U4105 ( .A1(n4353), .A2(sub_1_root_sub_0_root_u4_add_497_carry[8]), 
        .ZN(sub_1_root_sub_0_root_u4_add_497_carry[9]) );
  XNOR2_X1 U4106 ( .A(sub_1_root_sub_0_root_u4_add_497_carry[8]), .B(n4353), 
        .ZN(u4_ldz_dif_8_) );
  AND2_X1 U4107 ( .A1(n4281), .A2(u4_add_410_carry[7]), .ZN(
        u4_add_410_carry[8]) );
  XOR2_X1 U4108 ( .A(n4281), .B(u4_add_410_carry[7]), .Z(u4_div_shft2[7]) );
  AND2_X1 U4109 ( .A1(n4281), .A2(u4_add_411_carry[7]), .ZN(
        u4_add_411_carry[8]) );
  XOR2_X1 U4110 ( .A(n4281), .B(u4_add_411_carry[7]), .Z(u4_div_shft3_7_) );
  AND2_X1 U4111 ( .A1(u4_sub_412_carry[7]), .A2(n4348), .ZN(
        u4_sub_412_carry[8]) );
  XOR2_X1 U4112 ( .A(n4348), .B(u4_sub_412_carry[7]), .Z(u4_div_shft4[7]) );
  OR2_X1 U4113 ( .A1(n4281), .A2(sub_1_root_sub_0_root_u4_add_497_carry[7]), 
        .ZN(sub_1_root_sub_0_root_u4_add_497_carry[8]) );
  XNOR2_X1 U4114 ( .A(sub_1_root_sub_0_root_u4_add_497_carry[7]), .B(n4281), 
        .ZN(u4_ldz_dif_7_) );
  AND2_X1 U4115 ( .A1(exp_r[6]), .A2(u4_add_410_carry[6]), .ZN(
        u4_add_410_carry[7]) );
  XOR2_X1 U4116 ( .A(exp_r[6]), .B(u4_add_410_carry[6]), .Z(u4_div_shft2[6])
         );
  AND2_X1 U4117 ( .A1(n4290), .A2(u4_add_410_carry[5]), .ZN(
        u4_add_410_carry[6]) );
  XOR2_X1 U4118 ( .A(n4290), .B(u4_add_410_carry[5]), .Z(u4_div_shft2[5]) );
  AND2_X1 U4119 ( .A1(n4282), .A2(u4_add_410_carry[4]), .ZN(
        u4_add_410_carry[5]) );
  XOR2_X1 U4120 ( .A(n4282), .B(u4_add_410_carry[4]), .Z(u4_div_shft2[4]) );
  AND2_X1 U4121 ( .A1(n4655), .A2(u4_add_410_carry[3]), .ZN(
        u4_add_410_carry[4]) );
  XOR2_X1 U4122 ( .A(exp_r[3]), .B(u4_add_410_carry[3]), .Z(u4_div_shft2[3])
         );
  AND2_X1 U4123 ( .A1(n4315), .A2(exp_r[1]), .ZN(u4_add_410_carry[3]) );
  XOR2_X1 U4124 ( .A(n4315), .B(exp_r[1]), .Z(u4_div_shft2[2]) );
  AND2_X1 U4125 ( .A1(exp_r[6]), .A2(u4_add_411_carry[6]), .ZN(
        u4_add_411_carry[7]) );
  XOR2_X1 U4126 ( .A(exp_r[6]), .B(u4_add_411_carry[6]), .Z(u4_div_shft3_6_)
         );
  AND2_X1 U4127 ( .A1(n4290), .A2(u4_add_411_carry[5]), .ZN(
        u4_add_411_carry[6]) );
  XOR2_X1 U4128 ( .A(n4290), .B(u4_add_411_carry[5]), .Z(u4_div_shft3_5_) );
  AND2_X1 U4129 ( .A1(n4600), .A2(div_opa_ldz_r2[0]), .ZN(u4_add_411_carry[1])
         );
  XOR2_X1 U4130 ( .A(n4600), .B(div_opa_ldz_r2[0]), .Z(u4_div_shft3_0_) );
  XNOR2_X1 U4131 ( .A(u4_sub_409_carry[10]), .B(n4656), .ZN(u4_div_scht1a[10])
         );
  OR2_X1 U4132 ( .A1(n4289), .A2(u4_sub_409_carry[9]), .ZN(
        u4_sub_409_carry[10]) );
  XNOR2_X1 U4133 ( .A(u4_sub_409_carry[9]), .B(n4289), .ZN(u4_div_scht1a[9])
         );
  OR2_X1 U4134 ( .A1(n4353), .A2(u4_sub_409_carry[8]), .ZN(u4_sub_409_carry[9]) );
  XNOR2_X1 U4135 ( .A(u4_sub_409_carry[8]), .B(n4353), .ZN(u4_div_scht1a[8])
         );
  OR2_X1 U4136 ( .A1(n4281), .A2(u4_sub_409_carry[7]), .ZN(u4_sub_409_carry[8]) );
  XNOR2_X1 U4137 ( .A(u4_sub_409_carry[7]), .B(n4281), .ZN(u4_div_scht1a[7])
         );
  OR2_X1 U4138 ( .A1(exp_r[6]), .A2(u4_sub_409_carry[6]), .ZN(
        u4_sub_409_carry[7]) );
  XNOR2_X1 U4139 ( .A(u4_sub_409_carry[6]), .B(exp_r[6]), .ZN(u4_div_scht1a[6]) );
  OR2_X1 U4140 ( .A1(n4290), .A2(u4_sub_409_carry[5]), .ZN(u4_sub_409_carry[6]) );
  XNOR2_X1 U4141 ( .A(u4_sub_409_carry[5]), .B(n4290), .ZN(u4_div_scht1a[5])
         );
  OR2_X1 U4142 ( .A1(n4447), .A2(n4600), .ZN(u4_sub_409_carry[1]) );
  XNOR2_X1 U4143 ( .A(n4600), .B(n4447), .ZN(u4_div_scht1a[0]) );
  AND2_X1 U4144 ( .A1(u4_sub_412_carry[6]), .A2(n4317), .ZN(
        u4_sub_412_carry[7]) );
  XOR2_X1 U4145 ( .A(n4317), .B(u4_sub_412_carry[6]), .Z(u4_div_shft4[6]) );
  AND2_X1 U4146 ( .A1(u4_sub_412_carry[5]), .A2(n4347), .ZN(
        u4_sub_412_carry[6]) );
  XOR2_X1 U4147 ( .A(n4347), .B(u4_sub_412_carry[5]), .Z(u4_div_shft4[5]) );
  OR2_X1 U4148 ( .A1(n4349), .A2(div_opa_ldz_r2[0]), .ZN(u4_sub_412_carry[1])
         );
  XNOR2_X1 U4149 ( .A(div_opa_ldz_r2[0]), .B(n4349), .ZN(u4_div_shft4[0]) );
  XNOR2_X1 U4150 ( .A(n4656), .B(u4_sub_417_carry_10_), .ZN(u4_f2i_shft_10_)
         );
  OR2_X1 U4151 ( .A1(n4289), .A2(u4_sub_417_carry_9_), .ZN(
        u4_sub_417_carry_10_) );
  XNOR2_X1 U4152 ( .A(u4_sub_417_carry_9_), .B(n4289), .ZN(u4_f2i_shft_9_) );
  OR2_X1 U4153 ( .A1(n4353), .A2(u4_sub_417_carry_8_), .ZN(u4_sub_417_carry_9_) );
  XNOR2_X1 U4154 ( .A(u4_sub_417_carry_8_), .B(n4353), .ZN(u4_f2i_shft_8_) );
  OR2_X1 U4155 ( .A1(n4281), .A2(u4_sub_417_carry_7_), .ZN(u4_sub_417_carry_8_) );
  XNOR2_X1 U4156 ( .A(u4_sub_417_carry_7_), .B(n4281), .ZN(u4_f2i_shft_7_) );
  AND2_X1 U4157 ( .A1(u4_sub_417_carry_6_), .A2(exp_r[6]), .ZN(
        u4_sub_417_carry_7_) );
  XOR2_X1 U4158 ( .A(exp_r[6]), .B(u4_sub_417_carry_6_), .Z(u4_f2i_shft_6_) );
  AND2_X1 U4159 ( .A1(u4_sub_417_carry_5_), .A2(n4290), .ZN(
        u4_sub_417_carry_6_) );
  XOR2_X1 U4160 ( .A(n4290), .B(u4_sub_417_carry_5_), .Z(u4_f2i_shft_5_) );
  AND2_X1 U4161 ( .A1(u4_sub_417_carry_4_), .A2(n4282), .ZN(
        u4_sub_417_carry_5_) );
  XOR2_X1 U4162 ( .A(n4282), .B(u4_sub_417_carry_4_), .Z(u4_f2i_shft_4_) );
  AND2_X1 U4163 ( .A1(u4_sub_417_carry_3_), .A2(n4655), .ZN(
        u4_sub_417_carry_4_) );
  XOR2_X1 U4164 ( .A(n4655), .B(u4_sub_417_carry_3_), .Z(u4_f2i_shft_3_) );
  AND2_X1 U4165 ( .A1(u4_sub_417_carry_2_), .A2(n4315), .ZN(
        u4_sub_417_carry_3_) );
  XOR2_X1 U4166 ( .A(n4315), .B(u4_sub_417_carry_2_), .Z(u4_f2i_shft_2_) );
  OR2_X1 U4167 ( .A1(exp_r[1]), .A2(n4600), .ZN(u4_sub_417_carry_2_) );
  XNOR2_X1 U4168 ( .A(n4600), .B(exp_r[1]), .ZN(u4_f2i_shft_1_) );
  AND2_X1 U4169 ( .A1(u4_sub_481_carry[6]), .A2(n4663), .ZN(u4_N6142) );
  XOR2_X1 U4170 ( .A(n4663), .B(u4_sub_481_carry[6]), .Z(u4_N6141) );
  AND2_X1 U4171 ( .A1(u4_sub_481_carry[5]), .A2(n4664), .ZN(
        u4_sub_481_carry[6]) );
  XOR2_X1 U4172 ( .A(n4664), .B(u4_sub_481_carry[5]), .Z(u4_N6140) );
  OR2_X1 U4173 ( .A1(n4665), .A2(u4_sub_481_carry[4]), .ZN(u4_sub_481_carry[5]) );
  XNOR2_X1 U4174 ( .A(u4_sub_481_carry[4]), .B(n4665), .ZN(u4_N6139) );
  OR2_X1 U4175 ( .A1(n4714), .A2(u4_sub_481_carry[3]), .ZN(u4_sub_481_carry[4]) );
  XNOR2_X1 U4176 ( .A(u4_sub_481_carry[3]), .B(n4714), .ZN(u4_N6138) );
  OR2_X1 U4177 ( .A1(n4715), .A2(u4_sub_481_carry[2]), .ZN(u4_sub_481_carry[3]) );
  XNOR2_X1 U4178 ( .A(u4_sub_481_carry[2]), .B(n4715), .ZN(u4_N6137) );
  OR2_X1 U4179 ( .A1(n4666), .A2(u4_fi_ldz_mi1_0_), .ZN(u4_sub_481_carry[2])
         );
  XNOR2_X1 U4180 ( .A(u4_fi_ldz_mi1_0_), .B(n4666), .ZN(u4_N6136) );
  OR2_X1 U4181 ( .A1(exp_r[6]), .A2(sub_1_root_sub_0_root_u4_add_497_carry[6]), 
        .ZN(sub_1_root_sub_0_root_u4_add_497_carry[7]) );
  XNOR2_X1 U4182 ( .A(sub_1_root_sub_0_root_u4_add_497_carry[6]), .B(exp_r[6]), 
        .ZN(u4_ldz_dif_6_) );
  OR2_X1 U4183 ( .A1(n4290), .A2(sub_1_root_sub_0_root_u4_add_497_carry[5]), 
        .ZN(sub_1_root_sub_0_root_u4_add_497_carry[6]) );
  XNOR2_X1 U4184 ( .A(sub_1_root_sub_0_root_u4_add_497_carry[5]), .B(n4290), 
        .ZN(u4_ldz_dif_5_) );
  OR2_X1 U4185 ( .A1(n4447), .A2(n4600), .ZN(
        sub_1_root_sub_0_root_u4_add_497_carry[1]) );
  XNOR2_X1 U4186 ( .A(n4600), .B(n4447), .ZN(u4_ldz_dif_0_) );
  XOR2_X1 U4187 ( .A(n4663), .B(u4_sub_491_carry[6]), .Z(u4_fi_ldz_2a_6_) );
  OR2_X1 U4188 ( .A1(n4664), .A2(u4_sub_491_carry[5]), .ZN(u4_sub_491_carry[6]) );
  XNOR2_X1 U4189 ( .A(u4_sub_491_carry[5]), .B(n4664), .ZN(u4_fi_ldz_2a_5_) );
  OR2_X1 U4190 ( .A1(n4665), .A2(u4_sub_491_carry[4]), .ZN(u4_sub_491_carry[5]) );
  XNOR2_X1 U4191 ( .A(u4_sub_491_carry[4]), .B(n4665), .ZN(u4_fi_ldz_2a_4_) );
  AND2_X1 U4192 ( .A1(u4_sub_491_carry[3]), .A2(n4714), .ZN(
        u4_sub_491_carry[4]) );
  XOR2_X1 U4193 ( .A(n4714), .B(u4_sub_491_carry[3]), .Z(u4_fi_ldz_2a_3_) );
  OR2_X1 U4194 ( .A1(n4715), .A2(u4_sub_491_carry[2]), .ZN(u4_sub_491_carry[3]) );
  XNOR2_X1 U4195 ( .A(u4_sub_491_carry[2]), .B(n4715), .ZN(u4_fi_ldz_2a_2_) );
  AND2_X1 U4196 ( .A1(u4_fi_ldz_mi1_0_), .A2(n4666), .ZN(u4_sub_491_carry[2])
         );
  XOR2_X1 U4197 ( .A(n4666), .B(u4_fi_ldz_mi1_0_), .Z(u4_fi_ldz_2a_1_) );
  XNOR2_X1 U4198 ( .A(u2_gt_145_B_11_), .B(u2_sub_116_carry_11_), .ZN(u2_N53)
         );
  OR2_X1 U4199 ( .A1(u2_exp_tmp4_10_), .A2(u2_sub_116_carry_10_), .ZN(
        u2_sub_116_carry_11_) );
  XNOR2_X1 U4200 ( .A(u2_sub_116_carry_10_), .B(u2_exp_tmp4_10_), .ZN(u2_N52)
         );
  AND2_X1 U4201 ( .A1(u2_sub_116_carry_9_), .A2(u2_lt_135_A_9_), .ZN(
        u2_sub_116_carry_10_) );
  XOR2_X1 U4202 ( .A(u2_lt_135_A_9_), .B(u2_sub_116_carry_9_), .Z(u2_N51) );
  AND2_X1 U4203 ( .A1(u2_sub_116_carry_8_), .A2(u2_lt_135_A_8_), .ZN(
        u2_sub_116_carry_9_) );
  XOR2_X1 U4204 ( .A(u2_lt_135_A_8_), .B(u2_sub_116_carry_8_), .Z(u2_N50) );
  AND2_X1 U4205 ( .A1(u2_sub_116_carry_7_), .A2(u2_lt_135_A_7_), .ZN(
        u2_sub_116_carry_8_) );
  XOR2_X1 U4206 ( .A(u2_lt_135_A_7_), .B(u2_sub_116_carry_7_), .Z(u2_N49) );
  AND2_X1 U4207 ( .A1(u2_sub_116_carry_6_), .A2(u2_lt_135_A_6_), .ZN(
        u2_sub_116_carry_7_) );
  XOR2_X1 U4208 ( .A(u2_lt_135_A_6_), .B(u2_sub_116_carry_6_), .Z(u2_N48) );
  AND2_X1 U4209 ( .A1(u2_sub_116_carry_5_), .A2(u2_lt_135_A_5_), .ZN(
        u2_sub_116_carry_6_) );
  XOR2_X1 U4210 ( .A(u2_lt_135_A_5_), .B(u2_sub_116_carry_5_), .Z(u2_N47) );
  AND2_X1 U4211 ( .A1(u2_sub_116_carry_4_), .A2(u2_exp_tmp1_4_), .ZN(
        u2_sub_116_carry_5_) );
  XOR2_X1 U4212 ( .A(u2_exp_tmp1_4_), .B(u2_sub_116_carry_4_), .Z(u2_N46) );
  AND2_X1 U4213 ( .A1(u2_sub_116_carry_3_), .A2(u2_exp_tmp1_3_), .ZN(
        u2_sub_116_carry_4_) );
  XOR2_X1 U4214 ( .A(u2_exp_tmp1_3_), .B(u2_sub_116_carry_3_), .Z(u2_N45) );
  AND2_X1 U4215 ( .A1(u2_sub_116_carry_2_), .A2(u2_exp_tmp1_2_), .ZN(
        u2_sub_116_carry_3_) );
  XOR2_X1 U4216 ( .A(u2_exp_tmp1_2_), .B(u2_sub_116_carry_2_), .Z(u2_N44) );
  AND2_X1 U4217 ( .A1(u2_lt_135_A_0_), .A2(u2_exp_tmp1_1_), .ZN(
        u2_sub_116_carry_2_) );
  XOR2_X1 U4218 ( .A(u2_exp_tmp1_1_), .B(u2_lt_135_A_0_), .Z(u2_N43) );
  XOR2_X1 U4219 ( .A(u2_gt_145_B_11_), .B(u2_add_116_carry_11_), .Z(u2_N41) );
  AND2_X1 U4220 ( .A1(u2_add_116_carry_10_), .A2(u2_exp_tmp4_10_), .ZN(
        u2_add_116_carry_11_) );
  XOR2_X1 U4221 ( .A(u2_exp_tmp4_10_), .B(u2_add_116_carry_10_), .Z(u2_N40) );
  OR2_X1 U4222 ( .A1(u2_lt_135_A_9_), .A2(u2_add_116_carry_9_), .ZN(
        u2_add_116_carry_10_) );
  XNOR2_X1 U4223 ( .A(u2_add_116_carry_9_), .B(u2_lt_135_A_9_), .ZN(u2_N39) );
  OR2_X1 U4224 ( .A1(u2_lt_135_A_8_), .A2(u2_add_116_carry_8_), .ZN(
        u2_add_116_carry_9_) );
  XNOR2_X1 U4225 ( .A(u2_add_116_carry_8_), .B(u2_lt_135_A_8_), .ZN(u2_N38) );
  OR2_X1 U4226 ( .A1(u2_lt_135_A_7_), .A2(u2_add_116_carry_7_), .ZN(
        u2_add_116_carry_8_) );
  XNOR2_X1 U4227 ( .A(u2_add_116_carry_7_), .B(u2_lt_135_A_7_), .ZN(u2_N37) );
  OR2_X1 U4228 ( .A1(u2_lt_135_A_6_), .A2(u2_add_116_carry_6_), .ZN(
        u2_add_116_carry_7_) );
  XNOR2_X1 U4229 ( .A(u2_add_116_carry_6_), .B(u2_lt_135_A_6_), .ZN(u2_N36) );
  OR2_X1 U4230 ( .A1(u2_lt_135_A_5_), .A2(u2_add_116_carry_5_), .ZN(
        u2_add_116_carry_6_) );
  XNOR2_X1 U4231 ( .A(u2_add_116_carry_5_), .B(u2_lt_135_A_5_), .ZN(u2_N35) );
  OR2_X1 U4232 ( .A1(u2_exp_tmp1_4_), .A2(u2_add_116_carry_4_), .ZN(
        u2_add_116_carry_5_) );
  XNOR2_X1 U4233 ( .A(u2_add_116_carry_4_), .B(u2_exp_tmp1_4_), .ZN(u2_N34) );
  OR2_X1 U4234 ( .A1(u2_exp_tmp1_3_), .A2(u2_add_116_carry_3_), .ZN(
        u2_add_116_carry_4_) );
  XNOR2_X1 U4235 ( .A(u2_add_116_carry_3_), .B(u2_exp_tmp1_3_), .ZN(u2_N33) );
  OR2_X1 U4236 ( .A1(u2_exp_tmp1_2_), .A2(u2_add_116_carry_2_), .ZN(
        u2_add_116_carry_3_) );
  XNOR2_X1 U4237 ( .A(u2_add_116_carry_2_), .B(u2_exp_tmp1_2_), .ZN(u2_N32) );
  OR2_X1 U4238 ( .A1(u2_exp_tmp1_1_), .A2(u2_lt_135_A_0_), .ZN(
        u2_add_116_carry_2_) );
  XNOR2_X1 U4239 ( .A(u2_lt_135_A_0_), .B(u2_exp_tmp1_1_), .ZN(u2_N31) );
  INV_X4 U4240 ( .A(u4_fi_ldz_6_), .ZN(n4663) );
  INV_X4 U4241 ( .A(u4_fi_ldz_5_), .ZN(n4664) );
  INV_X4 U4242 ( .A(u4_fi_ldz_4_), .ZN(n4665) );
  INV_X4 U4243 ( .A(u4_fi_ldz_1_), .ZN(n4666) );
  INV_X4 U4244 ( .A(u2_exp_tmp1_1_), .ZN(u2_exp_tmp4_1_) );
  INV_X4 U4245 ( .A(u2_exp_tmp1_2_), .ZN(u2_exp_tmp4_2_) );
  INV_X4 U4246 ( .A(u2_exp_tmp1_3_), .ZN(u2_exp_tmp4_3_) );
  INV_X4 U4247 ( .A(u2_exp_tmp1_4_), .ZN(u2_exp_tmp4_4_) );
  NOR2_X1 U4248 ( .A1(u2_exp_tmp4_1_), .A2(n2800), .ZN(n4668) );
  NOR2_X1 U4249 ( .A1(n4677), .A2(u2_exp_tmp4_2_), .ZN(n4669) );
  NOR2_X1 U4250 ( .A1(n4678), .A2(u2_exp_tmp4_3_), .ZN(n4670) );
  NOR2_X1 U4251 ( .A1(n4378), .A2(n2799), .ZN(n4672) );
  NAND2_X1 U4252 ( .A1(n4672), .A2(u2_lt_135_A_6_), .ZN(n4673) );
  NOR2_X1 U4253 ( .A1(n4673), .A2(n2797), .ZN(n4675) );
  NAND2_X1 U4254 ( .A1(n4675), .A2(u2_lt_135_A_8_), .ZN(n4676) );
  NOR2_X1 U4255 ( .A1(n2795), .A2(n4676), .ZN(n4667) );
  XOR2_X1 U4256 ( .A(u2_exp_tmp4_10_), .B(n4667), .Z(u2_N75) );
  OAI21_X1 U4257 ( .B1(u2_lt_135_A_0_), .B2(u2_exp_tmp1_1_), .A(n4677), .ZN(
        u2_N66) );
  OAI21_X1 U4258 ( .B1(n4668), .B2(u2_exp_tmp1_2_), .A(n4678), .ZN(u2_N67) );
  OAI21_X1 U4259 ( .B1(n4669), .B2(u2_exp_tmp1_3_), .A(n4679), .ZN(u2_N68) );
  OAI21_X1 U4260 ( .B1(n4670), .B2(u2_exp_tmp1_4_), .A(n4378), .ZN(u2_N69) );
  AOI21_X1 U4261 ( .B1(n4378), .B2(n2799), .A(n4672), .ZN(n4671) );
  OAI21_X1 U4262 ( .B1(n4672), .B2(u2_lt_135_A_6_), .A(n4673), .ZN(u2_N71) );
  AOI21_X1 U4263 ( .B1(n4673), .B2(n2797), .A(n4675), .ZN(n4674) );
  OAI21_X1 U4264 ( .B1(n4675), .B2(u2_lt_135_A_8_), .A(n4676), .ZN(u2_N73) );
  XNOR2_X1 U4265 ( .A(n2795), .B(n4676), .ZN(u2_N74) );
  INV_X4 U4266 ( .A(n4668), .ZN(n4677) );
  INV_X4 U4267 ( .A(n4669), .ZN(n4678) );
  INV_X4 U4268 ( .A(n4670), .ZN(n4679) );
  INV_X4 U4269 ( .A(n4671), .ZN(u2_N70) );
  INV_X4 U4270 ( .A(n4674), .ZN(u2_N72) );
  NOR2_X1 U4271 ( .A1(exp_r[1]), .A2(n4600), .ZN(n4681) );
  NOR2_X1 U4272 ( .A1(u4_sub_417_carry_2_), .A2(n4315), .ZN(n4682) );
  NOR2_X1 U4273 ( .A1(n4689), .A2(n4655), .ZN(n4683) );
  NOR2_X1 U4274 ( .A1(n4690), .A2(n4282), .ZN(n4684) );
  NOR2_X1 U4275 ( .A1(n4691), .A2(n4290), .ZN(n4685) );
  NOR2_X1 U4276 ( .A1(n4354), .A2(n4281), .ZN(n4687) );
  NAND2_X1 U4277 ( .A1(n4687), .A2(n4439), .ZN(n4688) );
  NOR3_X1 U4278 ( .A1(n4352), .A2(n4289), .A3(n4688), .ZN(u4_exp_in_mi1_11_)
         );
  OAI21_X1 U4279 ( .B1(n4289), .B2(n4688), .A(n4352), .ZN(n4680) );
  NAND2_X1 U4280 ( .A1(n6460), .A2(n4680), .ZN(u4_exp_in_mi1_10_) );
  OAI21_X1 U4281 ( .B1(n4349), .B2(n4314), .A(u4_sub_417_carry_2_), .ZN(
        u4_exp_in_mi1_1_) );
  OAI21_X1 U4282 ( .B1(n4681), .B2(n4438), .A(n4689), .ZN(u4_exp_in_mi1_2_) );
  OAI21_X1 U4283 ( .B1(n4682), .B2(n4316), .A(n4690), .ZN(u4_exp_in_mi1_3_) );
  OAI21_X1 U4284 ( .B1(n4683), .B2(n4299), .A(n4691), .ZN(u4_exp_in_mi1_4_) );
  OAI21_X1 U4285 ( .B1(n4684), .B2(n4347), .A(n4692), .ZN(u4_exp_in_mi1_5_) );
  OAI21_X1 U4286 ( .B1(n4685), .B2(n4317), .A(n4354), .ZN(u4_exp_in_mi1_6_) );
  AOI21_X1 U4287 ( .B1(n4354), .B2(n4281), .A(n4687), .ZN(n4686) );
  OAI21_X1 U4288 ( .B1(n4687), .B2(n4439), .A(n4688), .ZN(u4_exp_in_mi1_8_) );
  XNOR2_X1 U4289 ( .A(n4289), .B(n4688), .ZN(u4_exp_in_mi1_9_) );
  INV_X4 U4290 ( .A(n4682), .ZN(n4689) );
  INV_X4 U4291 ( .A(n4683), .ZN(n4690) );
  INV_X4 U4292 ( .A(n4684), .ZN(n4691) );
  INV_X4 U4293 ( .A(n4685), .ZN(n4692) );
  INV_X4 U4294 ( .A(n4686), .ZN(u4_exp_in_mi1_7_) );
  NOR2_X1 U4295 ( .A1(u4_fi_ldz_1_), .A2(u4_fi_ldz_2a_0_), .ZN(n4694) );
  AOI21_X1 U4296 ( .B1(u4_fi_ldz_2a_0_), .B2(u4_fi_ldz_1_), .A(n4694), .ZN(
        n4693) );
  NAND2_X1 U4297 ( .A1(n4694), .A2(n4715), .ZN(n4695) );
  OAI21_X1 U4298 ( .B1(n4694), .B2(n4715), .A(n4695), .ZN(u4_fi_ldz_mi1_2_) );
  NOR2_X1 U4299 ( .A1(n4695), .A2(u4_fi_ldz_3_), .ZN(n4697) );
  AOI21_X1 U4300 ( .B1(n4695), .B2(u4_fi_ldz_3_), .A(n4697), .ZN(n4696) );
  NAND2_X1 U4301 ( .A1(n4697), .A2(n4665), .ZN(n4698) );
  OAI21_X1 U4302 ( .B1(n4697), .B2(n4665), .A(n4698), .ZN(u4_fi_ldz_mi1_4_) );
  XNOR2_X1 U4303 ( .A(u4_fi_ldz_5_), .B(n4698), .ZN(u4_fi_ldz_mi1_5_) );
  NOR2_X1 U4304 ( .A1(u4_fi_ldz_5_), .A2(n4698), .ZN(n4699) );
  XOR2_X1 U4305 ( .A(u4_fi_ldz_6_), .B(n4699), .Z(u4_fi_ldz_mi1_6_) );
  INV_X4 U4306 ( .A(u4_fi_ldz_2a_0_), .ZN(u4_fi_ldz_mi1_0_) );
  INV_X4 U4307 ( .A(n4693), .ZN(u4_fi_ldz_mi1_1_) );
  INV_X4 U4308 ( .A(n4696), .ZN(u4_fi_ldz_mi1_3_) );
  NOR2_X1 U4309 ( .A1(u4_exp_out1_1_), .A2(u4_exp_out1_0_), .ZN(n4701) );
  NOR2_X1 U4310 ( .A1(n4710), .A2(u4_sub_468_A_2_), .ZN(n4702) );
  NOR2_X1 U4311 ( .A1(n4712), .A2(u4_sub_468_A_3_), .ZN(n4703) );
  NOR2_X1 U4312 ( .A1(n4339), .A2(u4_sub_468_A_5_), .ZN(n4705) );
  NAND2_X1 U4313 ( .A1(n4705), .A2(n2418), .ZN(n4706) );
  NOR2_X1 U4314 ( .A1(n4706), .A2(u4_sub_468_A_7_), .ZN(n4708) );
  NAND2_X1 U4315 ( .A1(n4708), .A2(n2424), .ZN(n4709) );
  NOR2_X1 U4316 ( .A1(u4_sub_468_A_9_), .A2(n4709), .ZN(n4700) );
  XOR2_X1 U4317 ( .A(u4_sub_468_A_10_), .B(n4700), .Z(u4_exp_out1_mi1[10]) );
  OAI21_X1 U4318 ( .B1(u4_exp_out1_mi1[0]), .B2(n4711), .A(n4710), .ZN(
        u4_exp_out1_mi1[1]) );
  OAI21_X1 U4319 ( .B1(n4701), .B2(n2407), .A(n4712), .ZN(u4_exp_out1_mi1[2])
         );
  OAI21_X1 U4320 ( .B1(n4702), .B2(n2411), .A(n4713), .ZN(u4_exp_out1_mi1[3])
         );
  OAI21_X1 U4321 ( .B1(n4703), .B2(n2414), .A(n4339), .ZN(u4_exp_out1_mi1[4])
         );
  AOI21_X1 U4322 ( .B1(n4339), .B2(u4_sub_468_A_5_), .A(n4705), .ZN(n4704) );
  OAI21_X1 U4323 ( .B1(n4705), .B2(n2418), .A(n4706), .ZN(u4_exp_out1_mi1[6])
         );
  AOI21_X1 U4324 ( .B1(n4706), .B2(u4_sub_468_A_7_), .A(n4708), .ZN(n4707) );
  OAI21_X1 U4325 ( .B1(n4708), .B2(n2424), .A(n4709), .ZN(u4_exp_out1_mi1[8])
         );
  XNOR2_X1 U4326 ( .A(u4_sub_468_A_9_), .B(n4709), .ZN(u4_exp_out1_mi1[9]) );
  INV_X4 U4327 ( .A(u4_exp_out1_0_), .ZN(u4_exp_out1_mi1[0]) );
  INV_X4 U4328 ( .A(n4701), .ZN(n4710) );
  INV_X4 U4329 ( .A(u4_exp_out1_1_), .ZN(n4711) );
  INV_X4 U4330 ( .A(n4702), .ZN(n4712) );
  INV_X4 U4331 ( .A(n4703), .ZN(n4713) );
  INV_X4 U4332 ( .A(n4704), .ZN(u4_exp_out1_mi1[5]) );
  INV_X4 U4333 ( .A(n4707), .ZN(u4_exp_out1_mi1[7]) );
  INV_X4 U4334 ( .A(u4_fi_ldz_3_), .ZN(n4714) );
  INV_X4 U4335 ( .A(u4_fi_ldz_2_), .ZN(n4715) );
  INV_X1 U4336 ( .A(u4_exp_out_0_), .ZN(u4_exp_out_mi1[0]) );
  NOR2_X1 U4337 ( .A1(u4_exp_out_1_), .A2(u4_exp_out_0_), .ZN(n4719) );
  INV_X1 U4338 ( .A(n4719), .ZN(n4717) );
  NOR2_X1 U4339 ( .A1(n4717), .A2(u4_exp_out_2_), .ZN(n4721) );
  INV_X1 U4340 ( .A(n4721), .ZN(n4718) );
  NOR2_X1 U4341 ( .A1(n4718), .A2(u4_exp_out_3_), .ZN(n4722) );
  INV_X1 U4342 ( .A(n4722), .ZN(n4720) );
  NOR2_X1 U4343 ( .A1(n4337), .A2(u4_exp_out_5_), .ZN(n4724) );
  NAND2_X1 U4344 ( .A1(n4724), .A2(n2456), .ZN(n4725) );
  NOR2_X1 U4345 ( .A1(n4725), .A2(u4_exp_out_7_), .ZN(n4727) );
  NAND2_X1 U4346 ( .A1(n4727), .A2(n2450), .ZN(n4728) );
  NOR2_X1 U4347 ( .A1(u4_exp_out_9_), .A2(n4728), .ZN(n4716) );
  XOR2_X1 U4348 ( .A(u4_exp_out_10_), .B(n4716), .Z(u4_exp_out_mi1[10]) );
  OAI21_X1 U4349 ( .B1(u4_exp_out_mi1[0]), .B2(n2471), .A(n4717), .ZN(
        u4_exp_out_mi1[1]) );
  OAI21_X1 U4350 ( .B1(n4719), .B2(n2468), .A(n4718), .ZN(u4_exp_out_mi1[2])
         );
  OAI21_X1 U4351 ( .B1(n4721), .B2(n2465), .A(n4720), .ZN(u4_exp_out_mi1[3])
         );
  OAI21_X1 U4352 ( .B1(n4722), .B2(n2462), .A(n4337), .ZN(u4_exp_out_mi1[4])
         );
  AOI21_X1 U4353 ( .B1(n4337), .B2(u4_exp_out_5_), .A(n4724), .ZN(n4723) );
  INV_X1 U4354 ( .A(n4723), .ZN(u4_exp_out_mi1[5]) );
  OAI21_X1 U4355 ( .B1(n4724), .B2(n2456), .A(n4725), .ZN(u4_exp_out_mi1[6])
         );
  AOI21_X1 U4356 ( .B1(n4725), .B2(u4_exp_out_7_), .A(n4727), .ZN(n4726) );
  INV_X1 U4357 ( .A(n4726), .ZN(u4_exp_out_mi1[7]) );
  OAI21_X1 U4358 ( .B1(n4727), .B2(n2450), .A(n4728), .ZN(u4_exp_out_mi1[8])
         );
  XNOR2_X1 U4359 ( .A(u4_exp_out_9_), .B(n4728), .ZN(u4_exp_out_mi1[9]) );
  NAND2_X1 U4360 ( .A1(opb_r[54]), .A2(n4451), .ZN(n4745) );
  NAND2_X1 U4361 ( .A1(opb_r[59]), .A2(n4442), .ZN(n4747) );
  NAND2_X1 U4362 ( .A1(opb_r[60]), .A2(n4357), .ZN(n4748) );
  NAND2_X1 U4363 ( .A1(opb_r[57]), .A2(n4453), .ZN(n4742) );
  NAND2_X1 U4364 ( .A1(opb_r[58]), .A2(n4454), .ZN(n4740) );
  NAND2_X1 U4365 ( .A1(opb_r[55]), .A2(n4358), .ZN(n4741) );
  NAND2_X1 U4366 ( .A1(opb_r[56]), .A2(n4456), .ZN(n4744) );
  NOR2_X1 U4367 ( .A1(n4449), .A2(opb_r[52]), .ZN(n4730) );
  OAI21_X1 U4368 ( .B1(n4756), .B2(n4450), .A(opb_r[53]), .ZN(n4729) );
  OAI211_X1 U4369 ( .C1(opa_r[53]), .C2(n4730), .A(n4729), .B(n4745), .ZN(
        n4731) );
  OAI221_X1 U4370 ( .B1(opb_r[54]), .B2(n4451), .C1(opb_r[55]), .C2(n4358), 
        .A(n4731), .ZN(n4732) );
  NAND3_X1 U4371 ( .A1(n4741), .A2(n4744), .A3(n4732), .ZN(n4733) );
  OAI221_X1 U4372 ( .B1(opb_r[56]), .B2(n4456), .C1(opb_r[57]), .C2(n4453), 
        .A(n4733), .ZN(n4734) );
  NAND3_X1 U4373 ( .A1(n4742), .A2(n4740), .A3(n4734), .ZN(n4735) );
  OAI221_X1 U4374 ( .B1(opb_r[58]), .B2(n4454), .C1(opb_r[59]), .C2(n4442), 
        .A(n4735), .ZN(n4736) );
  NAND3_X1 U4375 ( .A1(n4747), .A2(n4748), .A3(n4736), .ZN(n4737) );
  OAI221_X1 U4376 ( .B1(opb_r[60]), .B2(n4357), .C1(opb_r[61]), .C2(n4448), 
        .A(n4737), .ZN(n4738) );
  NAND2_X1 U4377 ( .A1(opb_r[61]), .A2(n4448), .ZN(n4749) );
  OAI211_X1 U4378 ( .C1(opa_r[62]), .C2(n4755), .A(n4738), .B(n4749), .ZN(
        n4739) );
  AOI21_X1 U4379 ( .B1(n4755), .B2(opa_r[62]), .A(n4757), .ZN(n4754) );
  AND3_X1 U4380 ( .A1(n4742), .A2(n4741), .A3(n4740), .ZN(n4743) );
  NAND4_X1 U4381 ( .A1(n4745), .A2(n4754), .A3(n4744), .A4(n4743), .ZN(n4753)
         );
  AND2_X1 U4382 ( .A1(opb_r[52]), .A2(n4449), .ZN(n4746) );
  OAI22_X1 U4383 ( .A1(n4746), .A2(n4450), .B1(opb_r[53]), .B2(n4746), .ZN(
        n4751) );
  AND3_X1 U4384 ( .A1(n4749), .A2(n4748), .A3(n4747), .ZN(n4750) );
  OAI211_X1 U4385 ( .C1(opa_r[62]), .C2(n4755), .A(n4751), .B(n4750), .ZN(
        n4752) );
  NOR2_X1 U4386 ( .A1(n4753), .A2(n4752), .ZN(u1_N49) );
  INV_X4 U4387 ( .A(opb_r[62]), .ZN(n4755) );
  INV_X4 U4388 ( .A(n4730), .ZN(n4756) );
  INV_X4 U4389 ( .A(n4739), .ZN(n4757) );
  INV_X4 U4390 ( .A(n4754), .ZN(u1_expa_lt_expb) );
  NOR2_X1 U4391 ( .A1(u1_exp_diff_6_), .A2(u1_exp_diff_10_), .ZN(n4761) );
  OR3_X1 U4392 ( .A1(u1_exp_diff_2_), .A2(u1_exp_diff_1_), .A3(u1_exp_diff_0_), 
        .ZN(n4758) );
  NAND4_X1 U4393 ( .A1(u1_exp_diff_5_), .A2(u1_exp_diff_4_), .A3(
        u1_exp_diff_3_), .A4(n4758), .ZN(n4760) );
  NOR3_X1 U4394 ( .A1(u1_exp_diff_7_), .A2(u1_exp_diff_9_), .A3(u1_exp_diff_8_), .ZN(n4759) );
  NAND3_X1 U4395 ( .A1(n4761), .A2(n4760), .A3(n4759), .ZN(u1_exp_lt_27) );
  NOR2_X1 U4396 ( .A1(u4_div_shft3_6_), .A2(u4_div_shft3_10_), .ZN(n4764) );
  OAI211_X1 U4397 ( .C1(u4_div_shft3_2_), .C2(u4_div_shft3_3_), .A(
        u4_div_shft3_4_), .B(u4_div_shft3_5_), .ZN(n4763) );
  NOR3_X1 U4398 ( .A1(u4_div_shft3_7_), .A2(u4_div_shft3_9_), .A3(
        u4_div_shft3_8_), .ZN(n4762) );
  NAND3_X1 U4399 ( .A1(n4764), .A2(n4763), .A3(n4762), .ZN(u4_N5843) );
  NAND4_X1 U4400 ( .A1(u4_div_exp2_3_), .A2(u4_div_exp2_2_), .A3(
        u4_div_exp2_1_), .A4(u4_div_exp2_0_), .ZN(n4766) );
  NAND4_X1 U4401 ( .A1(u4_div_exp2_7_), .A2(u4_div_exp2_6_), .A3(
        u4_div_exp2_5_), .A4(u4_div_exp2_4_), .ZN(n4765) );
  NOR2_X1 U4402 ( .A1(n4766), .A2(n4765), .ZN(n4767) );
  OR4_X1 U4403 ( .A1(u4_div_exp2_10_), .A2(n4767), .A3(u4_div_exp2_9_), .A4(
        u4_div_exp2_8_), .ZN(u4_N6172) );
  NAND3_X1 U4404 ( .A1(u4_div_exp1_1_), .A2(u4_div_exp1_0_), .A3(
        u4_div_exp1_2_), .ZN(n4771) );
  NAND2_X1 U4405 ( .A1(u4_div_exp1_4_), .A2(u4_div_exp1_3_), .ZN(n4770) );
  NAND3_X1 U4406 ( .A1(u4_div_exp1_6_), .A2(u4_div_exp1_5_), .A3(
        u4_div_exp1_7_), .ZN(n4769) );
  NAND2_X1 U4407 ( .A1(u4_div_exp1_9_), .A2(u4_div_exp1_8_), .ZN(n4768) );
  NOR4_X1 U4408 ( .A1(n4771), .A2(n4770), .A3(n4769), .A4(n4768), .ZN(n4772)
         );
  NOR2_X1 U4409 ( .A1(u4_div_exp1_10_), .A2(n4772), .ZN(u4_N6194) );
  OAI211_X1 U4410 ( .C1(u4_ldz_all_3_), .C2(u4_ldz_all_2_), .A(u4_ldz_all_4_), 
        .B(u4_ldz_all_5_), .ZN(n4773) );
  NOR2_X1 U4411 ( .A1(u4_ldz_all_6_), .A2(n4774), .ZN(u4_N6286) );
  INV_X4 U4412 ( .A(n4773), .ZN(n4774) );
  OR3_X1 U4413 ( .A1(n4282), .A2(exp_r[3]), .A3(n4315), .ZN(n4775) );
  OR3_X1 U4414 ( .A1(exp_r[1]), .A2(n4600), .A3(n4775), .ZN(n4776) );
  AOI211_X1 U4415 ( .C1(n4290), .C2(n4776), .A(exp_r[6]), .B(n4352), .ZN(n4778) );
  NOR3_X1 U4416 ( .A1(n4281), .A2(n4289), .A3(n4353), .ZN(n4777) );
  NAND2_X1 U4417 ( .A1(n4778), .A2(n4777), .ZN(u4_N6284) );
  NAND4_X1 U4418 ( .A1(exp_r[3]), .A2(n4315), .A3(exp_r[1]), .A4(n4600), .ZN(
        n4780) );
  NAND3_X1 U4419 ( .A1(n4290), .A2(n4282), .A3(exp_r[6]), .ZN(n4779) );
  OAI21_X1 U4420 ( .B1(n4780), .B2(n4779), .A(n4440), .ZN(n4781) );
  NOR4_X1 U4421 ( .A1(n4781), .A2(n4281), .A3(n4289), .A4(n4353), .ZN(u4_N6283) );
  NOR2_X1 U4422 ( .A1(exp_r[6]), .A2(n4352), .ZN(n4783) );
  OAI211_X1 U4423 ( .C1(exp_r[3]), .C2(n4315), .A(n4282), .B(n4290), .ZN(n4782) );
  NAND2_X1 U4424 ( .A1(n4783), .A2(n4782), .ZN(n4784) );
  NOR4_X1 U4425 ( .A1(n4784), .A2(n4281), .A3(n4289), .A4(n4353), .ZN(u4_N6280) );
  NOR2_X1 U4426 ( .A1(n4290), .A2(n4352), .ZN(n4788) );
  AND3_X1 U4427 ( .A1(exp_r[1]), .A2(n4600), .A3(n4315), .ZN(n4785) );
  OAI21_X1 U4428 ( .B1(n4785), .B2(n4655), .A(n4282), .ZN(n4787) );
  NOR4_X1 U4429 ( .A1(n4289), .A2(n4353), .A3(n4281), .A4(exp_r[6]), .ZN(n4786) );
  NAND3_X1 U4430 ( .A1(n4788), .A2(n4787), .A3(n4786), .ZN(u4_N6278) );
  AND2_X1 U4431 ( .A1(u4_fi_ldz_2a_4_), .A2(u4_fi_ldz_2a_3_), .ZN(n4789) );
  OAI211_X1 U4432 ( .C1(u4_fi_ldz_2_), .C2(u4_fi_ldz_3_), .A(u4_fi_ldz_5_), 
        .B(u4_fi_ldz_4_), .ZN(n4790) );
  NAND2_X1 U4433 ( .A1(n4663), .A2(n4790), .ZN(u4_N6203) );
  OR4_X1 U4434 ( .A1(n4281), .A2(exp_r[6]), .A3(n4289), .A4(n4353), .ZN(n4797)
         );
  NOR2_X1 U4435 ( .A1(n4447), .A2(n4600), .ZN(n4791) );
  AOI21_X1 U4436 ( .B1(n4791), .B2(n4314), .A(div_opa_ldz_r2[1]), .ZN(n4792)
         );
  AOI221_X1 U4437 ( .B1(n4315), .B2(n4444), .C1(exp_r[1]), .C2(
        u4_sub_409_carry[1]), .A(n4792), .ZN(n4793) );
  AOI221_X1 U4438 ( .B1(div_opa_ldz_r2[3]), .B2(n4316), .C1(div_opa_ldz_r2[2]), 
        .C2(n4438), .A(n4793), .ZN(n4794) );
  AOI221_X1 U4439 ( .B1(n4282), .B2(n4445), .C1(n4655), .C2(n4443), .A(n4794), 
        .ZN(n4795) );
  AOI21_X1 U4440 ( .B1(div_opa_ldz_r2[4]), .B2(n4299), .A(n4795), .ZN(n4796)
         );
  NOR4_X1 U4441 ( .A1(n4797), .A2(n4796), .A3(n4290), .A4(n4352), .ZN(u4_N6171) );
  NAND3_X1 U4442 ( .A1(u2_exp_tmp1_1_), .A2(u2_lt_135_A_0_), .A3(
        u2_exp_tmp1_2_), .ZN(n4801) );
  NAND2_X1 U4443 ( .A1(u2_exp_tmp1_4_), .A2(u2_exp_tmp1_3_), .ZN(n4800) );
  NAND3_X1 U4444 ( .A1(u2_lt_135_A_6_), .A2(u2_lt_135_A_5_), .A3(
        u2_lt_135_A_7_), .ZN(n4799) );
  NAND2_X1 U4445 ( .A1(u2_lt_135_A_9_), .A2(u2_lt_135_A_8_), .ZN(n4798) );
  NOR4_X1 U4446 ( .A1(n4801), .A2(n4800), .A3(n4799), .A4(n4798), .ZN(n4802)
         );
  OAI21_X1 U4447 ( .B1(n4802), .B2(u2_exp_tmp4_10_), .A(u2_gt_145_B_11_), .ZN(
        n4803) );
  INV_X4 U4448 ( .A(n4803), .ZN(u2_N113) );
  NAND3_X1 U4449 ( .A1(u2_exp_tmp1_1_), .A2(u2_lt_135_A_0_), .A3(
        u2_exp_tmp1_2_), .ZN(n4807) );
  NAND2_X1 U4450 ( .A1(u2_exp_tmp1_4_), .A2(u2_exp_tmp1_3_), .ZN(n4806) );
  NAND3_X1 U4451 ( .A1(u2_lt_135_A_6_), .A2(u2_lt_135_A_5_), .A3(
        u2_lt_135_A_7_), .ZN(n4805) );
  NAND2_X1 U4452 ( .A1(u2_lt_135_A_9_), .A2(u2_lt_135_A_8_), .ZN(n4804) );
  NOR4_X1 U4453 ( .A1(n4807), .A2(n4806), .A3(n4805), .A4(n4804), .ZN(n4808)
         );
  NOR2_X1 U4454 ( .A1(u2_exp_tmp4_10_), .A2(n4808), .ZN(u2_N111) );
  OAI211_X1 U4455 ( .C1(u4_fi_ldz_3_), .C2(u4_fi_ldz_2_), .A(u4_fi_ldz_4_), 
        .B(u4_fi_ldz_5_), .ZN(n4809) );
  NOR2_X1 U4456 ( .A1(u4_fi_ldz_6_), .A2(n4810), .ZN(u4_N6279) );
  INV_X4 U4457 ( .A(n4809), .ZN(n4810) );
  OAI21_X1 U4458 ( .B1(u4_fi_ldz_2a_1_), .B2(u4_fi_ldz_2a_0_), .A(
        u4_fi_ldz_2a_2_), .ZN(n4811) );
  AOI21_X1 U4459 ( .B1(n4811), .B2(n4813), .A(n4814), .ZN(n4812) );
  INV_X4 U4460 ( .A(u4_fi_ldz_2a_3_), .ZN(n4813) );
  INV_X4 U4461 ( .A(u4_fi_ldz_2a_4_), .ZN(n4814) );
  NOR2_X1 U4462 ( .A1(exp_r[6]), .A2(n4290), .ZN(n4816) );
  NAND4_X1 U4463 ( .A1(exp_r[1]), .A2(n4315), .A3(n4282), .A4(n4655), .ZN(
        n4815) );
  AOI21_X1 U4464 ( .B1(n4816), .B2(n4815), .A(n4348), .ZN(n4817) );
  OR4_X1 U4465 ( .A1(n4352), .A2(n4817), .A3(n4289), .A4(n4353), .ZN(u4_N5837)
         );
  OAI211_X1 U4466 ( .C1(n4600), .C2(n4823), .A(exp_r[1]), .B(n4315), .ZN(n4821) );
  NAND2_X1 U4467 ( .A1(n4282), .A2(n4655), .ZN(n4820) );
  NAND3_X1 U4468 ( .A1(exp_r[6]), .A2(n4290), .A3(n4281), .ZN(n4819) );
  NAND2_X1 U4469 ( .A1(n4289), .A2(n4353), .ZN(n4818) );
  NOR4_X1 U4470 ( .A1(n4821), .A2(n4820), .A3(n4819), .A4(n4818), .ZN(n4822)
         );
  NOR2_X1 U4471 ( .A1(n4352), .A2(n4822), .ZN(u4_N5836) );
  INV_X4 U4472 ( .A(u4_N6410), .ZN(n4823) );
  NAND2_X2 U4473 ( .A1(u4_exp_f2i_1[116]), .A2(n2400), .ZN(n2429) );
  NAND2_X2 U4474 ( .A1(u4_exp_f2i_1[117]), .A2(n2400), .ZN(n2432) );
  NAND2_X2 U4475 ( .A1(u4_exp_f2i_1[115]), .A2(n2400), .ZN(n2425) );
  AOI22_X2 U4476 ( .A1(N343), .A2(n4552), .B1(N343), .B2(n4546), .ZN(n4249) );
  AOI22_X2 U4477 ( .A1(opa_r1[1]), .A2(n4553), .B1(N344), .B2(n4197), .ZN(
        n4248) );
  AOI22_X2 U4478 ( .A1(opa_r1[2]), .A2(n4553), .B1(N345), .B2(n4197), .ZN(
        n4247) );
  AOI22_X2 U4479 ( .A1(opa_r1[3]), .A2(n4553), .B1(N346), .B2(n4546), .ZN(
        n4246) );
  AOI22_X2 U4480 ( .A1(opa_r1[4]), .A2(n4553), .B1(N347), .B2(n4546), .ZN(
        n4245) );
  AOI22_X2 U4481 ( .A1(opa_r1[5]), .A2(n4552), .B1(N348), .B2(n4546), .ZN(
        n4244) );
  AOI22_X2 U4482 ( .A1(opa_r1[6]), .A2(n4553), .B1(N349), .B2(n4546), .ZN(
        n4243) );
  AOI22_X2 U4483 ( .A1(n4552), .A2(opa_r1[7]), .B1(N350), .B2(n4546), .ZN(
        n4242) );
  AOI22_X2 U4484 ( .A1(n4552), .A2(opa_r1[8]), .B1(N351), .B2(n4546), .ZN(
        n4241) );
  AOI22_X2 U4485 ( .A1(n4552), .A2(opa_r1[9]), .B1(N352), .B2(n4546), .ZN(
        n4240) );
  AOI22_X2 U4486 ( .A1(n4552), .A2(opa_r1[10]), .B1(N353), .B2(n4546), .ZN(
        n4239) );
  AOI22_X2 U4487 ( .A1(n4552), .A2(opa_r1[11]), .B1(N354), .B2(n4546), .ZN(
        n4238) );
  AOI22_X2 U4488 ( .A1(n4552), .A2(opa_r1[12]), .B1(N355), .B2(n4546), .ZN(
        n4237) );
  AOI22_X2 U4489 ( .A1(n4552), .A2(opa_r1[13]), .B1(N356), .B2(n4546), .ZN(
        n4236) );
  AOI22_X2 U4490 ( .A1(n4551), .A2(opa_r1[14]), .B1(N357), .B2(n4546), .ZN(
        n4235) );
  AOI22_X2 U4491 ( .A1(n4551), .A2(opa_r1[15]), .B1(N358), .B2(n4547), .ZN(
        n4234) );
  AOI22_X2 U4492 ( .A1(n4551), .A2(opa_r1[16]), .B1(N359), .B2(n4547), .ZN(
        n4233) );
  AOI22_X2 U4493 ( .A1(n4551), .A2(opa_r1[17]), .B1(N360), .B2(n4547), .ZN(
        n4232) );
  AOI22_X2 U4494 ( .A1(n4551), .A2(opa_r1[18]), .B1(N361), .B2(n4547), .ZN(
        n4231) );
  AOI22_X2 U4495 ( .A1(n4551), .A2(opa_r1[19]), .B1(N362), .B2(n4547), .ZN(
        n4230) );
  AOI22_X2 U4496 ( .A1(n4551), .A2(opa_r1[20]), .B1(N363), .B2(n4547), .ZN(
        n4229) );
  AOI22_X2 U4497 ( .A1(n4551), .A2(opa_r1[21]), .B1(N364), .B2(n4547), .ZN(
        n4228) );
  AOI22_X2 U4498 ( .A1(n4551), .A2(opa_r1[22]), .B1(N365), .B2(n4547), .ZN(
        n4227) );
  AOI22_X2 U4499 ( .A1(n4551), .A2(opa_r1[23]), .B1(N366), .B2(n4547), .ZN(
        n4226) );
  AOI22_X2 U4500 ( .A1(n4550), .A2(opa_r1[24]), .B1(N367), .B2(n4547), .ZN(
        n4225) );
  AOI22_X2 U4501 ( .A1(n4550), .A2(opa_r1[25]), .B1(N368), .B2(n4547), .ZN(
        n4224) );
  AOI22_X2 U4502 ( .A1(n4550), .A2(opa_r1[26]), .B1(N369), .B2(n4548), .ZN(
        n4223) );
  AOI22_X2 U4503 ( .A1(n4550), .A2(opa_r1[27]), .B1(N370), .B2(n4548), .ZN(
        n4222) );
  AOI22_X2 U4504 ( .A1(n4550), .A2(opa_r1[28]), .B1(N371), .B2(n4548), .ZN(
        n4221) );
  AOI22_X2 U4505 ( .A1(n4550), .A2(opa_r1[29]), .B1(N372), .B2(n4548), .ZN(
        n4220) );
  AOI22_X2 U4506 ( .A1(n4550), .A2(opa_r1[30]), .B1(N373), .B2(n4548), .ZN(
        n4219) );
  AOI22_X2 U4507 ( .A1(n4550), .A2(opa_r1[31]), .B1(N374), .B2(n4548), .ZN(
        n4218) );
  AOI22_X2 U4508 ( .A1(n4550), .A2(opa_r1[32]), .B1(N375), .B2(n4548), .ZN(
        n4217) );
  AOI22_X2 U4509 ( .A1(n4550), .A2(opa_r1[33]), .B1(N376), .B2(n4548), .ZN(
        n4216) );
  AOI22_X2 U4510 ( .A1(n4550), .A2(opa_r1[34]), .B1(N377), .B2(n4548), .ZN(
        n4215) );
  AOI22_X2 U4511 ( .A1(n4552), .A2(opa_r1[35]), .B1(N378), .B2(n4548), .ZN(
        n4214) );
  AOI22_X2 U4512 ( .A1(n4552), .A2(opa_r1[36]), .B1(N379), .B2(n4548), .ZN(
        n4213) );
  AOI22_X2 U4513 ( .A1(n4552), .A2(opa_r1[37]), .B1(N380), .B2(n4548), .ZN(
        n4212) );
  AOI22_X2 U4514 ( .A1(n4552), .A2(opa_r1[38]), .B1(N381), .B2(n4547), .ZN(
        n4211) );
  AOI22_X2 U4515 ( .A1(n4552), .A2(opa_r1[39]), .B1(N382), .B2(n4546), .ZN(
        n4210) );
  AOI22_X2 U4516 ( .A1(n4552), .A2(opa_r1[40]), .B1(N383), .B2(n4548), .ZN(
        n4209) );
  AOI22_X2 U4517 ( .A1(n4552), .A2(opa_r1[41]), .B1(N384), .B2(n4547), .ZN(
        n4208) );
  AOI22_X2 U4518 ( .A1(n4552), .A2(opa_r1[42]), .B1(N385), .B2(n4546), .ZN(
        n4207) );
  AOI22_X2 U4519 ( .A1(n4552), .A2(opa_r1[43]), .B1(N386), .B2(n4548), .ZN(
        n4206) );
  AOI22_X2 U4520 ( .A1(n4552), .A2(opa_r1[44]), .B1(N387), .B2(n4547), .ZN(
        n4205) );
  AOI22_X2 U4521 ( .A1(n4551), .A2(opa_r1[45]), .B1(N388), .B2(n4546), .ZN(
        n4204) );
  INV_X4 U4522 ( .A(n3504), .ZN(n5864) );
  INV_X4 U4523 ( .A(n2430), .ZN(n5865) );
  INV_X4 U4524 ( .A(n2427), .ZN(n5866) );
  INV_X4 U4525 ( .A(n2423), .ZN(n5867) );
  INV_X4 U4526 ( .A(n3512), .ZN(n5868) );
  INV_X4 U4527 ( .A(n3506), .ZN(n5869) );
  INV_X4 U4528 ( .A(n3509), .ZN(n5870) );
  INV_X4 U4529 ( .A(n2413), .ZN(n5871) );
  INV_X4 U4530 ( .A(n2410), .ZN(n5872) );
  INV_X4 U4531 ( .A(n2406), .ZN(n5873) );
  INV_X4 U4532 ( .A(N307), .ZN(n5874) );
  INV_X4 U4533 ( .A(N306), .ZN(n5875) );
  INV_X4 U4534 ( .A(n3192), .ZN(u6_N104) );
  INV_X4 U4535 ( .A(n3193), .ZN(u6_N103) );
  INV_X4 U4536 ( .A(n3194), .ZN(u6_N102) );
  INV_X4 U4537 ( .A(N302), .ZN(n5876) );
  INV_X4 U4538 ( .A(N301), .ZN(n5877) );
  INV_X4 U4539 ( .A(N300), .ZN(n5878) );
  INV_X4 U4540 ( .A(n3181), .ZN(u6_N98) );
  INV_X4 U4541 ( .A(N298), .ZN(n5879) );
  INV_X4 U4542 ( .A(N297), .ZN(n5880) );
  INV_X4 U4543 ( .A(n3182), .ZN(u6_N95) );
  INV_X4 U4544 ( .A(N295), .ZN(n5881) );
  INV_X4 U4545 ( .A(N294), .ZN(n5882) );
  INV_X4 U4546 ( .A(N293), .ZN(n5883) );
  INV_X4 U4547 ( .A(N292), .ZN(n5884) );
  INV_X4 U4548 ( .A(N291), .ZN(n5885) );
  INV_X4 U4549 ( .A(n3183), .ZN(u6_N89) );
  INV_X4 U4550 ( .A(n3184), .ZN(u6_N88) );
  INV_X4 U4551 ( .A(N288), .ZN(n5886) );
  INV_X4 U4552 ( .A(N287), .ZN(n5887) );
  INV_X4 U4553 ( .A(N286), .ZN(n5888) );
  INV_X4 U4554 ( .A(N285), .ZN(n5889) );
  INV_X4 U4555 ( .A(N284), .ZN(n5890) );
  INV_X4 U4556 ( .A(N283), .ZN(n5891) );
  INV_X4 U4557 ( .A(n3185), .ZN(u6_N81) );
  INV_X4 U4558 ( .A(N281), .ZN(n5892) );
  INV_X4 U4559 ( .A(n3186), .ZN(u6_N79) );
  INV_X4 U4560 ( .A(n3187), .ZN(u6_N78) );
  INV_X4 U4561 ( .A(N278), .ZN(n5893) );
  INV_X4 U4562 ( .A(N277), .ZN(n5894) );
  INV_X4 U4563 ( .A(N276), .ZN(n5895) );
  INV_X4 U4564 ( .A(n3188), .ZN(u6_N74) );
  INV_X4 U4565 ( .A(N274), .ZN(n5896) );
  INV_X4 U4566 ( .A(N273), .ZN(n5897) );
  INV_X4 U4567 ( .A(N272), .ZN(n5898) );
  INV_X4 U4568 ( .A(N271), .ZN(n5899) );
  INV_X4 U4569 ( .A(N270), .ZN(n5900) );
  INV_X4 U4570 ( .A(n3189), .ZN(u6_N68) );
  INV_X4 U4571 ( .A(N268), .ZN(n5901) );
  INV_X4 U4572 ( .A(N267), .ZN(n5902) );
  INV_X4 U4573 ( .A(N266), .ZN(n5903) );
  INV_X4 U4574 ( .A(N265), .ZN(n5904) );
  INV_X4 U4575 ( .A(N264), .ZN(n5905) );
  INV_X4 U4576 ( .A(N263), .ZN(n5906) );
  INV_X4 U4577 ( .A(N262), .ZN(n5907) );
  INV_X4 U4578 ( .A(N261), .ZN(n5908) );
  INV_X4 U4579 ( .A(n3190), .ZN(u6_N59) );
  INV_X4 U4580 ( .A(N259), .ZN(n5909) );
  INV_X4 U4581 ( .A(n3191), .ZN(u6_N57) );
  INV_X4 U4582 ( .A(N257), .ZN(n5910) );
  INV_X4 U4583 ( .A(N256), .ZN(n5911) );
  INV_X4 U4584 ( .A(n3783), .ZN(n5912) );
  INV_X4 U4585 ( .A(n4204), .ZN(n5913) );
  INV_X4 U4586 ( .A(n4205), .ZN(n5914) );
  INV_X4 U4587 ( .A(n4206), .ZN(n5915) );
  INV_X4 U4588 ( .A(n4207), .ZN(n5916) );
  INV_X4 U4589 ( .A(n4208), .ZN(n5917) );
  INV_X4 U4590 ( .A(n4209), .ZN(n5918) );
  INV_X4 U4591 ( .A(n4210), .ZN(n5919) );
  INV_X4 U4592 ( .A(n4211), .ZN(n5920) );
  INV_X4 U4593 ( .A(n4212), .ZN(n5921) );
  INV_X4 U4594 ( .A(n4213), .ZN(n5922) );
  INV_X4 U4595 ( .A(n4214), .ZN(n5923) );
  INV_X4 U4596 ( .A(n4215), .ZN(n5924) );
  INV_X4 U4597 ( .A(n4216), .ZN(n5925) );
  INV_X4 U4598 ( .A(n4217), .ZN(n5926) );
  INV_X4 U4599 ( .A(n4218), .ZN(n5927) );
  INV_X4 U4600 ( .A(n4219), .ZN(n5928) );
  INV_X4 U4601 ( .A(n4220), .ZN(n5929) );
  INV_X4 U4602 ( .A(n4221), .ZN(n5930) );
  INV_X4 U4603 ( .A(n4222), .ZN(n5931) );
  INV_X4 U4604 ( .A(n4223), .ZN(n5932) );
  INV_X4 U4605 ( .A(n4224), .ZN(n5933) );
  INV_X4 U4606 ( .A(n4225), .ZN(n5934) );
  INV_X4 U4607 ( .A(n4226), .ZN(n5935) );
  INV_X4 U4608 ( .A(n4227), .ZN(n5936) );
  INV_X4 U4609 ( .A(n4228), .ZN(n5937) );
  INV_X4 U4610 ( .A(n4229), .ZN(n5938) );
  INV_X4 U4611 ( .A(n4230), .ZN(n5939) );
  INV_X4 U4612 ( .A(n4231), .ZN(n5940) );
  INV_X4 U4613 ( .A(n4232), .ZN(n5941) );
  INV_X4 U4614 ( .A(n4233), .ZN(n5942) );
  INV_X4 U4615 ( .A(n4234), .ZN(n5943) );
  INV_X4 U4616 ( .A(n4235), .ZN(n5944) );
  INV_X4 U4617 ( .A(n4236), .ZN(n5945) );
  INV_X4 U4618 ( .A(n4237), .ZN(n5946) );
  INV_X4 U4619 ( .A(n4238), .ZN(n5947) );
  INV_X4 U4620 ( .A(n4239), .ZN(n5948) );
  INV_X4 U4621 ( .A(n4240), .ZN(n5949) );
  INV_X4 U4622 ( .A(n4241), .ZN(n5950) );
  INV_X4 U4623 ( .A(n4242), .ZN(n5951) );
  INV_X4 U4624 ( .A(n4243), .ZN(n5952) );
  INV_X4 U4625 ( .A(n4244), .ZN(n5953) );
  INV_X4 U4626 ( .A(n4245), .ZN(n5954) );
  INV_X4 U4627 ( .A(n4246), .ZN(n5955) );
  INV_X4 U4628 ( .A(n4247), .ZN(n5956) );
  INV_X4 U4629 ( .A(n4248), .ZN(n5957) );
  INV_X4 U4630 ( .A(N557), .ZN(n5958) );
  INV_X4 U4631 ( .A(N556), .ZN(n5959) );
  INV_X4 U4632 ( .A(N555), .ZN(n5960) );
  INV_X4 U4633 ( .A(N554), .ZN(n5961) );
  INV_X4 U4634 ( .A(N553), .ZN(n5962) );
  INV_X4 U4635 ( .A(N552), .ZN(n5963) );
  INV_X4 U4636 ( .A(N551), .ZN(n5964) );
  INV_X4 U4637 ( .A(N550), .ZN(n5965) );
  INV_X4 U4638 ( .A(N549), .ZN(n5966) );
  INV_X4 U4639 ( .A(N548), .ZN(n5967) );
  INV_X4 U4640 ( .A(N547), .ZN(n5968) );
  INV_X4 U4641 ( .A(N546), .ZN(n5969) );
  INV_X4 U4642 ( .A(N545), .ZN(n5970) );
  INV_X4 U4643 ( .A(N544), .ZN(n5971) );
  INV_X4 U4644 ( .A(N543), .ZN(n5972) );
  INV_X4 U4645 ( .A(N542), .ZN(n5973) );
  INV_X4 U4646 ( .A(N541), .ZN(n5974) );
  INV_X4 U4647 ( .A(N540), .ZN(n5975) );
  INV_X4 U4648 ( .A(N539), .ZN(n5976) );
  INV_X4 U4649 ( .A(N538), .ZN(n5977) );
  INV_X4 U4650 ( .A(N537), .ZN(n5978) );
  INV_X4 U4651 ( .A(N536), .ZN(n5979) );
  INV_X4 U4652 ( .A(N535), .ZN(n5980) );
  INV_X4 U4653 ( .A(N534), .ZN(n5981) );
  INV_X4 U4654 ( .A(N533), .ZN(n5982) );
  INV_X4 U4655 ( .A(N532), .ZN(n5983) );
  INV_X4 U4656 ( .A(N531), .ZN(n5984) );
  INV_X4 U4657 ( .A(N530), .ZN(n5985) );
  INV_X4 U4658 ( .A(N529), .ZN(n5986) );
  INV_X4 U4659 ( .A(N528), .ZN(n5987) );
  INV_X4 U4660 ( .A(N527), .ZN(n5988) );
  INV_X4 U4661 ( .A(N526), .ZN(n5989) );
  INV_X4 U4662 ( .A(N525), .ZN(n5990) );
  INV_X4 U4663 ( .A(N524), .ZN(n5991) );
  INV_X4 U4664 ( .A(N523), .ZN(n5992) );
  INV_X4 U4665 ( .A(N522), .ZN(n5993) );
  INV_X4 U4666 ( .A(N521), .ZN(n5994) );
  INV_X4 U4667 ( .A(N520), .ZN(n5995) );
  INV_X4 U4668 ( .A(N519), .ZN(n5996) );
  INV_X4 U4669 ( .A(N518), .ZN(n5997) );
  INV_X4 U4670 ( .A(N517), .ZN(n5998) );
  INV_X4 U4671 ( .A(N516), .ZN(n5999) );
  INV_X4 U4672 ( .A(N515), .ZN(n6000) );
  INV_X4 U4673 ( .A(N514), .ZN(n6001) );
  INV_X4 U4674 ( .A(N513), .ZN(n6002) );
  INV_X4 U4675 ( .A(N512), .ZN(n6003) );
  INV_X4 U4676 ( .A(N511), .ZN(n6004) );
  INV_X4 U4677 ( .A(N510), .ZN(n6005) );
  INV_X4 U4678 ( .A(N509), .ZN(n6006) );
  INV_X4 U4679 ( .A(N508), .ZN(n6007) );
  INV_X4 U4680 ( .A(N507), .ZN(n6008) );
  INV_X4 U4681 ( .A(N506), .ZN(n6009) );
  INV_X4 U4682 ( .A(N505), .ZN(n6010) );
  INV_X4 U4683 ( .A(N504), .ZN(n6011) );
  INV_X4 U4684 ( .A(N503), .ZN(n6012) );
  INV_X4 U4685 ( .A(N502), .ZN(n6013) );
  INV_X4 U4686 ( .A(N501), .ZN(n6014) );
  INV_X4 U4687 ( .A(u2_exp_ovf_d_1_), .ZN(n6015) );
  INV_X4 U4688 ( .A(n2784), .ZN(u2_gt_145_B_11_) );
  INV_X4 U4689 ( .A(n2804), .ZN(n6016) );
  INV_X4 U4690 ( .A(u2_N16), .ZN(n6017) );
  INV_X4 U4691 ( .A(n2785), .ZN(n6018) );
  INV_X4 U4692 ( .A(n2795), .ZN(u2_lt_135_A_9_) );
  INV_X4 U4693 ( .A(n2786), .ZN(n6019) );
  INV_X4 U4694 ( .A(n2796), .ZN(u2_lt_135_A_8_) );
  INV_X4 U4695 ( .A(n2787), .ZN(n6020) );
  INV_X4 U4696 ( .A(n2797), .ZN(u2_lt_135_A_7_) );
  INV_X4 U4697 ( .A(n2788), .ZN(n6021) );
  INV_X4 U4698 ( .A(n2798), .ZN(u2_lt_135_A_6_) );
  INV_X4 U4699 ( .A(n2789), .ZN(n6022) );
  INV_X4 U4700 ( .A(n2799), .ZN(u2_lt_135_A_5_) );
  INV_X4 U4701 ( .A(n2790), .ZN(n6023) );
  INV_X4 U4702 ( .A(u2_N10), .ZN(n6024) );
  INV_X4 U4703 ( .A(n2791), .ZN(n6025) );
  INV_X4 U4704 ( .A(u2_N9), .ZN(n6026) );
  INV_X4 U4705 ( .A(n2792), .ZN(n6027) );
  INV_X4 U4706 ( .A(u2_N8), .ZN(n6028) );
  INV_X4 U4707 ( .A(n2793), .ZN(n6029) );
  INV_X4 U4708 ( .A(u2_N7), .ZN(n6030) );
  INV_X4 U4709 ( .A(n2794), .ZN(n6031) );
  INV_X4 U4710 ( .A(u2_N28), .ZN(n6032) );
  INV_X4 U4711 ( .A(u2_N22), .ZN(n6033) );
  INV_X4 U4712 ( .A(u2_N21), .ZN(n6034) );
  INV_X4 U4713 ( .A(u2_N20), .ZN(n6035) );
  INV_X4 U4714 ( .A(u2_N19), .ZN(n6036) );
  INV_X4 U4715 ( .A(n3292), .ZN(n6037) );
  INV_X4 U4716 ( .A(n3119), .ZN(n6038) );
  INV_X4 U4717 ( .A(n3120), .ZN(n6039) );
  INV_X4 U4718 ( .A(n3121), .ZN(n6040) );
  INV_X4 U4719 ( .A(n3122), .ZN(n6041) );
  INV_X4 U4720 ( .A(n3123), .ZN(n6042) );
  INV_X4 U4721 ( .A(n3124), .ZN(n6043) );
  INV_X4 U4722 ( .A(n3126), .ZN(n6044) );
  INV_X4 U4723 ( .A(n3127), .ZN(n6045) );
  INV_X4 U4724 ( .A(n3128), .ZN(n6046) );
  INV_X4 U4725 ( .A(n3129), .ZN(n6047) );
  INV_X4 U4726 ( .A(n3130), .ZN(n6048) );
  INV_X4 U4727 ( .A(n3131), .ZN(n6049) );
  INV_X4 U4728 ( .A(n3132), .ZN(n6050) );
  INV_X4 U4729 ( .A(n3133), .ZN(n6051) );
  INV_X4 U4730 ( .A(n3134), .ZN(n6052) );
  INV_X4 U4731 ( .A(n3135), .ZN(n6053) );
  INV_X4 U4732 ( .A(n3137), .ZN(n6054) );
  INV_X4 U4733 ( .A(n3138), .ZN(n6055) );
  INV_X4 U4734 ( .A(n3139), .ZN(n6056) );
  INV_X4 U4735 ( .A(n3140), .ZN(n6057) );
  INV_X4 U4736 ( .A(n3141), .ZN(n6058) );
  INV_X4 U4737 ( .A(n3142), .ZN(n6059) );
  INV_X4 U4738 ( .A(n3143), .ZN(n6060) );
  INV_X4 U4739 ( .A(n3144), .ZN(n6061) );
  INV_X4 U4740 ( .A(n3145), .ZN(n6062) );
  INV_X4 U4741 ( .A(n3146), .ZN(n6063) );
  INV_X4 U4742 ( .A(n3148), .ZN(n6064) );
  INV_X4 U4743 ( .A(n3149), .ZN(n6065) );
  INV_X4 U4744 ( .A(n3150), .ZN(n6066) );
  INV_X4 U4745 ( .A(n3151), .ZN(n6067) );
  INV_X4 U4746 ( .A(n3152), .ZN(n6068) );
  INV_X4 U4747 ( .A(n3153), .ZN(n6069) );
  INV_X4 U4748 ( .A(n3154), .ZN(n6070) );
  INV_X4 U4749 ( .A(n3155), .ZN(n6071) );
  INV_X4 U4750 ( .A(n3156), .ZN(n6072) );
  INV_X4 U4751 ( .A(n3157), .ZN(n6073) );
  INV_X4 U4752 ( .A(n3159), .ZN(n6074) );
  INV_X4 U4753 ( .A(n3160), .ZN(n6075) );
  INV_X4 U4754 ( .A(n3161), .ZN(n6076) );
  INV_X4 U4755 ( .A(n3162), .ZN(n6077) );
  INV_X4 U4756 ( .A(n3163), .ZN(n6078) );
  INV_X4 U4757 ( .A(n3164), .ZN(n6079) );
  INV_X4 U4758 ( .A(n3165), .ZN(n6080) );
  INV_X4 U4759 ( .A(n3166), .ZN(n6081) );
  INV_X4 U4760 ( .A(n3167), .ZN(n6082) );
  INV_X4 U4761 ( .A(n3168), .ZN(n6083) );
  INV_X4 U4762 ( .A(n3114), .ZN(n6084) );
  INV_X4 U4763 ( .A(n3115), .ZN(n6085) );
  INV_X4 U4764 ( .A(n3116), .ZN(n6086) );
  INV_X4 U4765 ( .A(n3117), .ZN(n6087) );
  INV_X4 U4766 ( .A(n3118), .ZN(n6088) );
  INV_X4 U4767 ( .A(n3125), .ZN(n6089) );
  INV_X4 U4768 ( .A(n3136), .ZN(n6090) );
  INV_X4 U4769 ( .A(n3147), .ZN(n6091) );
  INV_X4 U4770 ( .A(n3158), .ZN(n6092) );
  INV_X4 U4771 ( .A(n3169), .ZN(n6093) );
  INV_X4 U4772 ( .A(n3545), .ZN(n6094) );
  INV_X4 U4773 ( .A(n2438), .ZN(n6095) );
  INV_X4 U4774 ( .A(u4_exp_next_mi_11_), .ZN(n6096) );
  INV_X4 U4775 ( .A(n2431), .ZN(u4_sub_468_A_10_) );
  INV_X4 U4776 ( .A(n2428), .ZN(u4_sub_468_A_9_) );
  INV_X4 U4777 ( .A(n2420), .ZN(u4_sub_468_A_7_) );
  INV_X4 U4778 ( .A(n2416), .ZN(u4_sub_468_A_5_) );
  INV_X4 U4779 ( .A(n2414), .ZN(u4_sub_468_A_4_) );
  INV_X4 U4780 ( .A(n2411), .ZN(u4_sub_468_A_3_) );
  INV_X4 U4781 ( .A(n2407), .ZN(u4_sub_468_A_2_) );
  INV_X4 U4782 ( .A(u4_exp_next_mi_1_), .ZN(n6097) );
  INV_X4 U4783 ( .A(u4_exp_next_mi_0_), .ZN(n6098) );
  INV_X4 U4784 ( .A(u1_N232), .ZN(n6099) );
  INV_X4 U4785 ( .A(n2836), .ZN(n6100) );
  INV_X4 U4786 ( .A(n2838), .ZN(n6101) );
  INV_X4 U4787 ( .A(n2840), .ZN(n6102) );
  INV_X4 U4788 ( .A(n2842), .ZN(n6103) );
  INV_X4 U4789 ( .A(n2844), .ZN(n6104) );
  INV_X4 U4790 ( .A(n2846), .ZN(n6105) );
  INV_X4 U4791 ( .A(n2848), .ZN(n6106) );
  INV_X4 U4792 ( .A(n2850), .ZN(n6107) );
  INV_X4 U4793 ( .A(n2852), .ZN(n6108) );
  INV_X4 U4794 ( .A(n2854), .ZN(n6109) );
  INV_X4 U4795 ( .A(n2856), .ZN(n6110) );
  INV_X4 U4796 ( .A(n2858), .ZN(n6111) );
  INV_X4 U4797 ( .A(n2860), .ZN(n6112) );
  INV_X4 U4798 ( .A(n2862), .ZN(n6113) );
  INV_X4 U4799 ( .A(n2864), .ZN(n6114) );
  INV_X4 U4800 ( .A(n2866), .ZN(n6115) );
  INV_X4 U4801 ( .A(n2868), .ZN(n6116) );
  INV_X4 U4802 ( .A(n2870), .ZN(n6117) );
  INV_X4 U4803 ( .A(n2872), .ZN(n6118) );
  INV_X4 U4804 ( .A(n2874), .ZN(n6119) );
  INV_X4 U4805 ( .A(n2876), .ZN(n6120) );
  INV_X4 U4806 ( .A(n2878), .ZN(n6121) );
  INV_X4 U4807 ( .A(n2880), .ZN(n6122) );
  INV_X4 U4808 ( .A(n2882), .ZN(n6123) );
  INV_X4 U4809 ( .A(n2884), .ZN(n6124) );
  INV_X4 U4810 ( .A(n2886), .ZN(n6125) );
  INV_X4 U4811 ( .A(n2888), .ZN(n6126) );
  INV_X4 U4812 ( .A(n2890), .ZN(n6127) );
  INV_X4 U4813 ( .A(n2892), .ZN(n6128) );
  INV_X4 U4814 ( .A(n2894), .ZN(n6129) );
  INV_X4 U4815 ( .A(n2896), .ZN(n6130) );
  INV_X4 U4816 ( .A(n2898), .ZN(n6131) );
  INV_X4 U4817 ( .A(n2900), .ZN(n6132) );
  INV_X4 U4818 ( .A(n2904), .ZN(n6133) );
  INV_X4 U4819 ( .A(n2906), .ZN(n6134) );
  INV_X4 U4820 ( .A(n2908), .ZN(n6135) );
  INV_X4 U4821 ( .A(n2910), .ZN(n6136) );
  INV_X4 U4822 ( .A(n2912), .ZN(n6137) );
  INV_X4 U4823 ( .A(n2914), .ZN(n6138) );
  INV_X4 U4824 ( .A(n2916), .ZN(n6139) );
  INV_X4 U4825 ( .A(n2918), .ZN(n6140) );
  INV_X4 U4826 ( .A(n2920), .ZN(n6141) );
  INV_X4 U4827 ( .A(n2922), .ZN(n6142) );
  INV_X4 U4828 ( .A(n2926), .ZN(n6143) );
  INV_X4 U4829 ( .A(n2928), .ZN(n6144) );
  INV_X4 U4830 ( .A(n2930), .ZN(n6145) );
  INV_X4 U4831 ( .A(n2932), .ZN(n6146) );
  INV_X4 U4832 ( .A(n2934), .ZN(n6147) );
  INV_X4 U4833 ( .A(n2936), .ZN(n6148) );
  INV_X4 U4834 ( .A(n2938), .ZN(n6149) );
  INV_X4 U4835 ( .A(n2940), .ZN(n6150) );
  INV_X4 U4836 ( .A(n2942), .ZN(n6151) );
  INV_X4 U4837 ( .A(n2944), .ZN(n6152) );
  INV_X4 U4838 ( .A(n2837), .ZN(n6153) );
  INV_X4 U4839 ( .A(n2839), .ZN(n6154) );
  INV_X4 U4840 ( .A(n2841), .ZN(n6155) );
  INV_X4 U4841 ( .A(n2843), .ZN(n6156) );
  INV_X4 U4842 ( .A(n2845), .ZN(n6157) );
  INV_X4 U4843 ( .A(n2847), .ZN(n6158) );
  INV_X4 U4844 ( .A(n2849), .ZN(n6159) );
  INV_X4 U4845 ( .A(n2851), .ZN(n6160) );
  INV_X4 U4846 ( .A(n2853), .ZN(n6161) );
  INV_X4 U4847 ( .A(n2855), .ZN(n6162) );
  INV_X4 U4848 ( .A(n2857), .ZN(n6163) );
  INV_X4 U4849 ( .A(n2859), .ZN(n6164) );
  INV_X4 U4850 ( .A(n2861), .ZN(n6165) );
  INV_X4 U4851 ( .A(n2863), .ZN(n6166) );
  INV_X4 U4852 ( .A(n2865), .ZN(n6167) );
  INV_X4 U4853 ( .A(n2867), .ZN(n6168) );
  INV_X4 U4854 ( .A(n2869), .ZN(n6169) );
  INV_X4 U4855 ( .A(n2871), .ZN(n6170) );
  INV_X4 U4856 ( .A(n2873), .ZN(n6171) );
  INV_X4 U4857 ( .A(n2875), .ZN(n6172) );
  INV_X4 U4858 ( .A(n2877), .ZN(n6173) );
  INV_X4 U4859 ( .A(n2879), .ZN(n6174) );
  INV_X4 U4860 ( .A(n2881), .ZN(n6175) );
  INV_X4 U4861 ( .A(n2883), .ZN(n6176) );
  INV_X4 U4862 ( .A(n2885), .ZN(n6177) );
  INV_X4 U4863 ( .A(n2887), .ZN(n6178) );
  INV_X4 U4864 ( .A(n2889), .ZN(n6179) );
  INV_X4 U4865 ( .A(n2891), .ZN(n6180) );
  INV_X4 U4866 ( .A(n2893), .ZN(n6181) );
  INV_X4 U4867 ( .A(n2895), .ZN(n6182) );
  INV_X4 U4868 ( .A(n2897), .ZN(n6183) );
  INV_X4 U4869 ( .A(n2899), .ZN(n6184) );
  INV_X4 U4870 ( .A(n2901), .ZN(n6185) );
  INV_X4 U4871 ( .A(n2903), .ZN(n6186) );
  INV_X4 U4872 ( .A(n2905), .ZN(n6187) );
  INV_X4 U4873 ( .A(n2907), .ZN(n6188) );
  INV_X4 U4874 ( .A(n2909), .ZN(n6189) );
  INV_X4 U4875 ( .A(n2911), .ZN(n6190) );
  INV_X4 U4876 ( .A(n2913), .ZN(n6191) );
  INV_X4 U4877 ( .A(n2915), .ZN(n6192) );
  INV_X4 U4878 ( .A(n2917), .ZN(n6193) );
  INV_X4 U4879 ( .A(n2919), .ZN(n6194) );
  INV_X4 U4880 ( .A(n2921), .ZN(n6195) );
  INV_X4 U4881 ( .A(n2923), .ZN(n6196) );
  INV_X4 U4882 ( .A(n2925), .ZN(n6197) );
  INV_X4 U4883 ( .A(n2927), .ZN(n6198) );
  INV_X4 U4884 ( .A(n2929), .ZN(n6199) );
  INV_X4 U4885 ( .A(n2931), .ZN(n6200) );
  INV_X4 U4886 ( .A(n2933), .ZN(n6201) );
  INV_X4 U4887 ( .A(n2935), .ZN(n6202) );
  INV_X4 U4888 ( .A(n2937), .ZN(n6203) );
  INV_X4 U4889 ( .A(n2939), .ZN(n6204) );
  INV_X4 U4890 ( .A(n2941), .ZN(n6205) );
  INV_X4 U4891 ( .A(n2943), .ZN(n6206) );
  INV_X4 U4892 ( .A(n2945), .ZN(n6207) );
  INV_X4 U4893 ( .A(n2947), .ZN(n6208) );
  INV_X4 U4894 ( .A(n2946), .ZN(n6209) );
  INV_X4 U4895 ( .A(n2924), .ZN(n6210) );
  INV_X4 U4896 ( .A(n2902), .ZN(n6211) );
  INV_X4 U4897 ( .A(n2968), .ZN(n6212) );
  INV_X4 U4898 ( .A(n2980), .ZN(n6213) );
  INV_X4 U4899 ( .A(n2975), .ZN(n6214) );
  INV_X4 U4900 ( .A(n2974), .ZN(n6215) );
  INV_X4 U4901 ( .A(n2960), .ZN(n6216) );
  INV_X4 U4902 ( .A(n3003), .ZN(n6217) );
  INV_X4 U4903 ( .A(n2961), .ZN(n6218) );
  INV_X4 U4904 ( .A(n2966), .ZN(n6219) );
  INV_X4 U4905 ( .A(n2958), .ZN(n6220) );
  INV_X4 U4906 ( .A(n2953), .ZN(n6221) );
  INV_X4 U4907 ( .A(n2995), .ZN(n6222) );
  INV_X4 U4908 ( .A(u1_exp_lt_27), .ZN(n6223) );
  INV_X4 U4909 ( .A(n3001), .ZN(n6224) );
  INV_X4 U4910 ( .A(n3012), .ZN(n6225) );
  INV_X4 U4911 ( .A(n3004), .ZN(n6226) );
  INV_X4 U4912 ( .A(n3048), .ZN(n6227) );
  INV_X4 U4913 ( .A(n3049), .ZN(n6228) );
  INV_X4 U4914 ( .A(n3035), .ZN(n6229) );
  INV_X4 U4915 ( .A(n3034), .ZN(n6230) );
  INV_X4 U4916 ( .A(n3033), .ZN(n6231) );
  INV_X4 U4917 ( .A(n3032), .ZN(n6232) );
  INV_X4 U4918 ( .A(n3053), .ZN(n6233) );
  INV_X4 U4919 ( .A(n3013), .ZN(n6234) );
  INV_X4 U4920 ( .A(n3054), .ZN(n6235) );
  INV_X4 U4921 ( .A(n3055), .ZN(n6236) );
  INV_X4 U4922 ( .A(n3014), .ZN(n6237) );
  INV_X4 U4923 ( .A(n3056), .ZN(n6238) );
  INV_X4 U4924 ( .A(n3015), .ZN(n6239) );
  INV_X4 U4925 ( .A(n3016), .ZN(n6240) );
  INV_X4 U4926 ( .A(n3017), .ZN(n6241) );
  INV_X4 U4927 ( .A(n3018), .ZN(n6242) );
  INV_X4 U4928 ( .A(n3057), .ZN(n6243) );
  INV_X4 U4929 ( .A(n3019), .ZN(n6244) );
  INV_X4 U4930 ( .A(n3020), .ZN(n6245) );
  INV_X4 U4931 ( .A(n3021), .ZN(n6246) );
  INV_X4 U4932 ( .A(n3058), .ZN(n6247) );
  INV_X4 U4933 ( .A(n3022), .ZN(n6248) );
  INV_X4 U4934 ( .A(n3023), .ZN(n6249) );
  INV_X4 U4935 ( .A(n3038), .ZN(n6250) );
  INV_X4 U4936 ( .A(n3024), .ZN(n6251) );
  INV_X4 U4937 ( .A(n3025), .ZN(n6252) );
  INV_X4 U4938 ( .A(n3026), .ZN(n6253) );
  INV_X4 U4939 ( .A(n3037), .ZN(n6254) );
  INV_X4 U4940 ( .A(n3039), .ZN(n6255) );
  INV_X4 U4941 ( .A(n3042), .ZN(n6256) );
  INV_X4 U4942 ( .A(n3041), .ZN(n6257) );
  INV_X4 U4943 ( .A(n3043), .ZN(n6258) );
  INV_X4 U4944 ( .A(n3046), .ZN(n6259) );
  INV_X4 U4945 ( .A(n3045), .ZN(n6260) );
  INV_X4 U4946 ( .A(n3047), .ZN(n6261) );
  INV_X4 U4947 ( .A(u1_exp_large_10_), .ZN(n6262) );
  INV_X4 U4948 ( .A(n3050), .ZN(n6263) );
  INV_X4 U4949 ( .A(n3051), .ZN(n6264) );
  INV_X4 U4950 ( .A(u1_exp_large_7_), .ZN(n6265) );
  INV_X4 U4951 ( .A(u1_exp_large_6_), .ZN(n6266) );
  INV_X4 U4952 ( .A(u1_exp_large_5_), .ZN(n6267) );
  INV_X4 U4953 ( .A(u1_exp_large_4_), .ZN(n6268) );
  INV_X4 U4954 ( .A(u1_exp_large_3_), .ZN(n6269) );
  INV_X4 U4955 ( .A(u1_exp_large_2_), .ZN(n6270) );
  INV_X4 U4956 ( .A(u1_exp_large_1_), .ZN(n6271) );
  INV_X4 U4957 ( .A(u1_exp_large_0_), .ZN(n6272) );
  INV_X4 U4958 ( .A(n4266), .ZN(n6273) );
  INV_X4 U4959 ( .A(n2783), .ZN(n6274) );
  INV_X4 U4960 ( .A(u1_N46), .ZN(n6275) );
  INV_X4 U4961 ( .A(n3075), .ZN(n6276) );
  INV_X4 U4962 ( .A(n3242), .ZN(n6277) );
  INV_X4 U4963 ( .A(n3227), .ZN(n6278) );
  INV_X4 U4964 ( .A(n3260), .ZN(n6279) );
  INV_X4 U4965 ( .A(n3208), .ZN(n6280) );
  INV_X4 U4966 ( .A(n3272), .ZN(n6281) );
  INV_X4 U4967 ( .A(n3209), .ZN(n6282) );
  INV_X4 U4968 ( .A(n3229), .ZN(n6283) );
  INV_X4 U4969 ( .A(n3220), .ZN(n6284) );
  INV_X4 U4970 ( .A(n3236), .ZN(n6285) );
  INV_X4 U4971 ( .A(n3266), .ZN(n6286) );
  INV_X4 U4972 ( .A(n3284), .ZN(n6287) );
  INV_X4 U4973 ( .A(n3204), .ZN(n6288) );
  INV_X4 U4974 ( .A(n3268), .ZN(n6289) );
  INV_X4 U4975 ( .A(n3239), .ZN(n6290) );
  INV_X4 U4976 ( .A(n3259), .ZN(n6291) );
  INV_X4 U4977 ( .A(n3207), .ZN(n6292) );
  INV_X4 U4978 ( .A(n3226), .ZN(n6293) );
  INV_X4 U4979 ( .A(n3218), .ZN(n6294) );
  INV_X4 U4980 ( .A(n3240), .ZN(n6295) );
  INV_X4 U4981 ( .A(n3237), .ZN(n6296) );
  INV_X4 U4982 ( .A(n3092), .ZN(n6297) );
  INV_X4 U4983 ( .A(n3283), .ZN(n6298) );
  INV_X4 U4984 ( .A(n3289), .ZN(n6299) );
  INV_X4 U4985 ( .A(n3246), .ZN(n6300) );
  INV_X4 U4986 ( .A(n3090), .ZN(n6301) );
  INV_X4 U4987 ( .A(n3222), .ZN(n6302) );
  INV_X4 U4988 ( .A(u6_N52), .ZN(n6303) );
  INV_X4 U4989 ( .A(n3074), .ZN(n6304) );
  INV_X4 U4990 ( .A(n3741), .ZN(n6305) );
  INV_X4 U4991 ( .A(n3737), .ZN(n6306) );
  INV_X4 U4992 ( .A(n2435), .ZN(n6307) );
  INV_X4 U4993 ( .A(u4_N5836), .ZN(n6308) );
  INV_X4 U4994 ( .A(n3548), .ZN(n6309) );
  INV_X4 U4995 ( .A(n3619), .ZN(n6310) );
  INV_X4 U4996 ( .A(n4249), .ZN(n6311) );
  INV_X4 U4997 ( .A(n4190), .ZN(n6313) );
  INV_X4 U4998 ( .A(n3343), .ZN(n6314) );
  INV_X4 U4999 ( .A(n2507), .ZN(n6316) );
  INV_X4 U5000 ( .A(n3297), .ZN(n6317) );
  INV_X4 U5001 ( .A(u4_N6203), .ZN(n6318) );
  INV_X4 U5002 ( .A(n2699), .ZN(n6319) );
  INV_X4 U5003 ( .A(n2651), .ZN(n6320) );
  INV_X4 U5004 ( .A(n2688), .ZN(n6321) );
  INV_X4 U5005 ( .A(n2572), .ZN(n6322) );
  INV_X4 U5006 ( .A(n2690), .ZN(n6323) );
  INV_X4 U5007 ( .A(n2617), .ZN(n6324) );
  INV_X4 U5008 ( .A(n2642), .ZN(n6325) );
  INV_X4 U5009 ( .A(n2679), .ZN(n6326) );
  INV_X4 U5010 ( .A(n2632), .ZN(n6327) );
  INV_X4 U5011 ( .A(n2555), .ZN(n6328) );
  INV_X4 U5012 ( .A(n2600), .ZN(n6329) );
  INV_X4 U5013 ( .A(n2613), .ZN(n6330) );
  INV_X4 U5014 ( .A(n2615), .ZN(n6331) );
  INV_X4 U5015 ( .A(n2639), .ZN(n6332) );
  INV_X4 U5016 ( .A(n2585), .ZN(n6333) );
  INV_X4 U5017 ( .A(n2562), .ZN(n6334) );
  INV_X4 U5018 ( .A(n2647), .ZN(n6335) );
  INV_X4 U5019 ( .A(n2671), .ZN(n6336) );
  INV_X4 U5020 ( .A(n2422), .ZN(n6337) );
  INV_X4 U5021 ( .A(n2598), .ZN(n6338) );
  INV_X4 U5022 ( .A(n2439), .ZN(n6339) );
  INV_X4 U5023 ( .A(n2447), .ZN(n6340) );
  INV_X4 U5024 ( .A(n3311), .ZN(n6341) );
  INV_X4 U5025 ( .A(n2433), .ZN(n6343) );
  INV_X4 U5026 ( .A(n3879), .ZN(n6344) );
  INV_X4 U5027 ( .A(n2724), .ZN(n6345) );
  INV_X4 U5028 ( .A(n3873), .ZN(n6346) );
  INV_X4 U5029 ( .A(n2763), .ZN(n6347) );
  INV_X4 U5030 ( .A(n3171), .ZN(n6348) );
  INV_X4 U5031 ( .A(n2751), .ZN(n6349) );
  INV_X4 U5032 ( .A(n2767), .ZN(n6350) );
  INV_X4 U5033 ( .A(n2683), .ZN(n6351) );
  INV_X4 U5034 ( .A(n2599), .ZN(n6352) );
  INV_X4 U5035 ( .A(fract_denorm[91]), .ZN(n6353) );
  INV_X4 U5036 ( .A(fract_denorm[92]), .ZN(n6354) );
  INV_X4 U5037 ( .A(fract_denorm[94]), .ZN(n6355) );
  INV_X4 U5038 ( .A(fract_denorm[96]), .ZN(n6356) );
  INV_X4 U5039 ( .A(n2738), .ZN(n6357) );
  INV_X4 U5040 ( .A(fract_denorm[97]), .ZN(n6358) );
  INV_X4 U5041 ( .A(fract_denorm[90]), .ZN(n6359) );
  INV_X4 U5042 ( .A(fract_denorm[99]), .ZN(n6360) );
  INV_X4 U5043 ( .A(fract_denorm[103]), .ZN(n6361) );
  INV_X4 U5044 ( .A(fract_denorm[104]), .ZN(n6362) );
  INV_X4 U5045 ( .A(fract_denorm[101]), .ZN(n6363) );
  INV_X4 U5046 ( .A(fract_denorm[100]), .ZN(n6364) );
  INV_X4 U5047 ( .A(fract_denorm[98]), .ZN(n6365) );
  INV_X4 U5048 ( .A(n2771), .ZN(n6366) );
  INV_X4 U5049 ( .A(n2711), .ZN(n6367) );
  INV_X4 U5050 ( .A(n4097), .ZN(n6368) );
  INV_X4 U5051 ( .A(n3912), .ZN(n6369) );
  INV_X4 U5052 ( .A(fract_denorm[54]), .ZN(n6370) );
  INV_X4 U5053 ( .A(fract_denorm[56]), .ZN(n6371) );
  INV_X4 U5054 ( .A(n2750), .ZN(n6372) );
  INV_X4 U5055 ( .A(fract_denorm[57]), .ZN(n6373) );
  INV_X4 U5056 ( .A(fract_denorm[84]), .ZN(n6374) );
  INV_X4 U5057 ( .A(n2760), .ZN(n6375) );
  INV_X4 U5058 ( .A(fract_denorm[86]), .ZN(n6376) );
  INV_X4 U5059 ( .A(fract_denorm[88]), .ZN(n6377) );
  INV_X4 U5060 ( .A(n2749), .ZN(n6378) );
  INV_X4 U5061 ( .A(fract_denorm[89]), .ZN(n6379) );
  INV_X4 U5062 ( .A(n2560), .ZN(n6380) );
  INV_X4 U5063 ( .A(fract_denorm[76]), .ZN(n6381) );
  INV_X4 U5064 ( .A(n2728), .ZN(n6382) );
  INV_X4 U5065 ( .A(fract_denorm[78]), .ZN(n6383) );
  INV_X4 U5066 ( .A(fract_denorm[80]), .ZN(n6384) );
  INV_X4 U5067 ( .A(n2736), .ZN(n6385) );
  INV_X4 U5068 ( .A(fract_denorm[79]), .ZN(n6386) );
  INV_X4 U5069 ( .A(fract_denorm[59]), .ZN(n6387) );
  INV_X4 U5070 ( .A(n2705), .ZN(n6388) );
  INV_X4 U5071 ( .A(fract_denorm[62]), .ZN(n6389) );
  INV_X4 U5072 ( .A(fract_denorm[64]), .ZN(n6390) );
  INV_X4 U5073 ( .A(n2735), .ZN(n6391) );
  INV_X4 U5074 ( .A(fract_denorm[63]), .ZN(n6392) );
  INV_X4 U5075 ( .A(n2646), .ZN(n6393) );
  INV_X4 U5076 ( .A(fract_denorm[68]), .ZN(n6394) );
  INV_X4 U5077 ( .A(fract_denorm[69]), .ZN(n6395) );
  INV_X4 U5078 ( .A(n2759), .ZN(n6396) );
  INV_X4 U5079 ( .A(fract_denorm[72]), .ZN(n6397) );
  INV_X4 U5080 ( .A(n2661), .ZN(n6398) );
  INV_X4 U5081 ( .A(fract_denorm[71]), .ZN(n6399) );
  INV_X4 U5082 ( .A(fract_denorm[52]), .ZN(n6400) );
  INV_X4 U5083 ( .A(fract_denorm[58]), .ZN(n6401) );
  INV_X4 U5084 ( .A(fract_denorm[82]), .ZN(n6402) );
  INV_X4 U5085 ( .A(fract_denorm[51]), .ZN(n6403) );
  INV_X4 U5086 ( .A(fract_denorm[50]), .ZN(n6404) );
  INV_X4 U5087 ( .A(n3173), .ZN(n6405) );
  INV_X4 U5088 ( .A(n2729), .ZN(n6406) );
  INV_X4 U5089 ( .A(n3172), .ZN(n6407) );
  INV_X4 U5090 ( .A(n2737), .ZN(n6408) );
  INV_X4 U5091 ( .A(n2744), .ZN(n6409) );
  INV_X4 U5092 ( .A(n4095), .ZN(n6410) );
  INV_X4 U5093 ( .A(n3180), .ZN(n6411) );
  INV_X4 U5094 ( .A(n2561), .ZN(n6412) );
  INV_X4 U5095 ( .A(n2731), .ZN(n6413) );
  INV_X4 U5096 ( .A(n3179), .ZN(n6414) );
  INV_X4 U5097 ( .A(n2740), .ZN(n6415) );
  INV_X4 U5098 ( .A(n2745), .ZN(n6416) );
  INV_X4 U5099 ( .A(n2593), .ZN(n6417) );
  INV_X4 U5100 ( .A(n4008), .ZN(n6418) );
  INV_X4 U5101 ( .A(n3178), .ZN(n6419) );
  INV_X4 U5102 ( .A(n2762), .ZN(n6420) );
  INV_X4 U5103 ( .A(n3177), .ZN(n6421) );
  INV_X4 U5104 ( .A(n2753), .ZN(n6422) );
  INV_X4 U5105 ( .A(n2769), .ZN(n6423) );
  INV_X4 U5106 ( .A(n2685), .ZN(n6424) );
  INV_X4 U5107 ( .A(n4000), .ZN(n6425) );
  INV_X4 U5108 ( .A(n3176), .ZN(n6426) );
  INV_X4 U5109 ( .A(n2730), .ZN(n6427) );
  INV_X4 U5110 ( .A(n3175), .ZN(n6428) );
  INV_X4 U5111 ( .A(n2739), .ZN(n6429) );
  INV_X4 U5112 ( .A(n2681), .ZN(n6430) );
  INV_X4 U5113 ( .A(n2722), .ZN(n6431) );
  INV_X4 U5114 ( .A(n3992), .ZN(n6432) );
  INV_X4 U5115 ( .A(n2758), .ZN(n6433) );
  INV_X4 U5116 ( .A(n2696), .ZN(n6434) );
  INV_X4 U5117 ( .A(n3174), .ZN(n6435) );
  INV_X4 U5118 ( .A(n2752), .ZN(n6436) );
  INV_X4 U5119 ( .A(n2680), .ZN(n6437) );
  INV_X4 U5120 ( .A(n2768), .ZN(n6438) );
  INV_X4 U5121 ( .A(n3984), .ZN(n6439) );
  INV_X4 U5122 ( .A(n2633), .ZN(n6440) );
  INV_X4 U5123 ( .A(n2605), .ZN(n6441) );
  INV_X4 U5124 ( .A(n2636), .ZN(n6442) );
  INV_X4 U5125 ( .A(n3876), .ZN(n6443) );
  INV_X4 U5126 ( .A(n2718), .ZN(n6444) );
  INV_X4 U5127 ( .A(n2770), .ZN(n6445) );
  INV_X4 U5128 ( .A(n3877), .ZN(n6446) );
  INV_X4 U5129 ( .A(n3488), .ZN(n6447) );
  INV_X4 U5130 ( .A(n3913), .ZN(n6448) );
  INV_X4 U5131 ( .A(n3459), .ZN(n6449) );
  INV_X4 U5132 ( .A(n3068), .ZN(n6450) );
  INV_X4 U5133 ( .A(n3069), .ZN(n6451) );
  INV_X4 U5134 ( .A(n3070), .ZN(n6452) );
  INV_X4 U5135 ( .A(n3071), .ZN(n6453) );
  INV_X4 U5136 ( .A(n3306), .ZN(n6454) );
  INV_X4 U5137 ( .A(n3565), .ZN(n6455) );
  INV_X4 U5138 ( .A(n3457), .ZN(n6456) );
  INV_X4 U5139 ( .A(n3314), .ZN(n6457) );
  INV_X4 U5140 ( .A(n3303), .ZN(n6458) );
  INV_X4 U5141 ( .A(n3454), .ZN(n6459) );
  INV_X4 U5142 ( .A(u4_exp_in_mi1_11_), .ZN(n6460) );
  INV_X4 U5143 ( .A(u4_exp_in_pl1_4_), .ZN(n6461) );
  INV_X4 U5144 ( .A(u4_exp_in_pl1_3_), .ZN(n6462) );
  INV_X4 U5145 ( .A(u4_exp_in_pl1_2_), .ZN(n6463) );
  INV_X4 U5146 ( .A(u4_exp_in_pl1_1_), .ZN(n6464) );
  INV_X4 U5147 ( .A(n2514), .ZN(n6465) );
  INV_X4 U5148 ( .A(n3787), .ZN(n6466) );
  INV_X4 U5149 ( .A(u4_N5837), .ZN(n6467) );
  INV_X4 U5150 ( .A(n3965), .ZN(n6468) );
  INV_X4 u4_sub_473_U23 ( .A(u4_fi_ldz_mi1_0_), .ZN(u4_sub_473_n14) );
  INV_X4 u4_sub_473_U22 ( .A(u4_fi_ldz_mi1_1_), .ZN(u4_sub_473_n13) );
  INV_X4 u4_sub_473_U21 ( .A(u4_fi_ldz_mi1_6_), .ZN(u4_sub_473_n12) );
  INV_X4 u4_sub_473_U20 ( .A(u4_fi_ldz_mi1_5_), .ZN(u4_sub_473_n11) );
  INV_X4 u4_sub_473_U19 ( .A(u4_fi_ldz_mi1_4_), .ZN(u4_sub_473_n10) );
  INV_X4 u4_sub_473_U18 ( .A(u4_fi_ldz_mi1_3_), .ZN(u4_sub_473_n9) );
  INV_X4 u4_sub_473_U17 ( .A(u4_fi_ldz_mi1_2_), .ZN(u4_sub_473_n8) );
  INV_X4 u4_sub_473_U16 ( .A(n4600), .ZN(u4_sub_473_n7) );
  XNOR2_X2 u4_sub_473_U15 ( .A(u4_sub_473_n14), .B(n4600), .ZN(
        u4_exp_fix_divb[0]) );
  NAND2_X2 u4_sub_473_U14 ( .A1(u4_fi_ldz_mi1_0_), .A2(u4_sub_473_n7), .ZN(
        u4_sub_473_carry_1_) );
  INV_X4 u4_sub_473_U13 ( .A(u4_sub_473_carry_9_), .ZN(u4_sub_473_n6) );
  INV_X4 u4_sub_473_U12 ( .A(n4289), .ZN(u4_sub_473_n5) );
  XNOR2_X2 u4_sub_473_U11 ( .A(n4289), .B(u4_sub_473_carry_9_), .ZN(
        u4_exp_fix_divb[9]) );
  NAND2_X2 u4_sub_473_U10 ( .A1(u4_sub_473_n5), .A2(u4_sub_473_n6), .ZN(
        u4_sub_473_carry_10_) );
  INV_X4 u4_sub_473_U9 ( .A(u4_sub_473_carry_8_), .ZN(u4_sub_473_n4) );
  INV_X4 u4_sub_473_U8 ( .A(n4353), .ZN(u4_sub_473_n3) );
  XNOR2_X2 u4_sub_473_U7 ( .A(n4353), .B(u4_sub_473_carry_8_), .ZN(
        u4_exp_fix_divb[8]) );
  NAND2_X2 u4_sub_473_U6 ( .A1(u4_sub_473_n3), .A2(u4_sub_473_n4), .ZN(
        u4_sub_473_carry_9_) );
  INV_X4 u4_sub_473_U5 ( .A(u4_sub_473_carry_7_), .ZN(u4_sub_473_n2) );
  INV_X4 u4_sub_473_U4 ( .A(n4281), .ZN(u4_sub_473_n1) );
  XNOR2_X2 u4_sub_473_U3 ( .A(n4281), .B(u4_sub_473_carry_7_), .ZN(
        u4_exp_fix_divb[7]) );
  NAND2_X2 u4_sub_473_U2 ( .A1(u4_sub_473_n1), .A2(u4_sub_473_n2), .ZN(
        u4_sub_473_carry_8_) );
  XNOR2_X2 u4_sub_473_U1 ( .A(n4656), .B(u4_sub_473_carry_10_), .ZN(
        u4_exp_fix_divb[10]) );
  FA_X1 u4_sub_473_U2_1 ( .A(exp_r[1]), .B(u4_sub_473_n13), .CI(
        u4_sub_473_carry_1_), .CO(u4_sub_473_carry_2_), .S(u4_exp_fix_divb[1])
         );
  FA_X1 u4_sub_473_U2_2 ( .A(n4315), .B(u4_sub_473_n8), .CI(
        u4_sub_473_carry_2_), .CO(u4_sub_473_carry_3_), .S(u4_exp_fix_divb[2])
         );
  FA_X1 u4_sub_473_U2_3 ( .A(n4655), .B(u4_sub_473_n9), .CI(
        u4_sub_473_carry_3_), .CO(u4_sub_473_carry_4_), .S(u4_exp_fix_divb[3])
         );
  FA_X1 u4_sub_473_U2_4 ( .A(n4282), .B(u4_sub_473_n10), .CI(
        u4_sub_473_carry_4_), .CO(u4_sub_473_carry_5_), .S(u4_exp_fix_divb[4])
         );
  FA_X1 u4_sub_473_U2_5 ( .A(n4290), .B(u4_sub_473_n11), .CI(
        u4_sub_473_carry_5_), .CO(u4_sub_473_carry_6_), .S(u4_exp_fix_divb[5])
         );
  FA_X1 u4_sub_473_U2_6 ( .A(exp_r[6]), .B(u4_sub_473_n12), .CI(
        u4_sub_473_carry_6_), .CO(u4_sub_473_carry_7_), .S(u4_exp_fix_divb[6])
         );
  INV_X4 u4_sub_472_U23 ( .A(u4_fi_ldz_mi1_0_), .ZN(u4_sub_472_n14) );
  INV_X4 u4_sub_472_U22 ( .A(u4_fi_ldz_mi22[1]), .ZN(u4_sub_472_n13) );
  INV_X4 u4_sub_472_U21 ( .A(u4_fi_ldz_mi22[2]), .ZN(u4_sub_472_n12) );
  INV_X4 u4_sub_472_U20 ( .A(u4_fi_ldz_mi22[3]), .ZN(u4_sub_472_n11) );
  INV_X4 u4_sub_472_U19 ( .A(u4_fi_ldz_mi22[4]), .ZN(u4_sub_472_n10) );
  INV_X4 u4_sub_472_U18 ( .A(u4_fi_ldz_mi22[5]), .ZN(u4_sub_472_n9) );
  INV_X4 u4_sub_472_U17 ( .A(u4_fi_ldz_mi22[6]), .ZN(u4_sub_472_n8) );
  INV_X4 u4_sub_472_U16 ( .A(n4600), .ZN(u4_sub_472_n7) );
  XNOR2_X2 u4_sub_472_U15 ( .A(u4_sub_472_n14), .B(n4600), .ZN(
        u4_exp_fix_diva[0]) );
  NAND2_X2 u4_sub_472_U14 ( .A1(u4_fi_ldz_mi1_0_), .A2(u4_sub_472_n7), .ZN(
        u4_sub_472_carry_1_) );
  INV_X4 u4_sub_472_U13 ( .A(u4_sub_472_carry_9_), .ZN(u4_sub_472_n6) );
  INV_X4 u4_sub_472_U12 ( .A(n4289), .ZN(u4_sub_472_n5) );
  XNOR2_X2 u4_sub_472_U11 ( .A(n4289), .B(u4_sub_472_carry_9_), .ZN(
        u4_exp_fix_diva[9]) );
  NAND2_X2 u4_sub_472_U10 ( .A1(u4_sub_472_n5), .A2(u4_sub_472_n6), .ZN(
        u4_sub_472_carry_10_) );
  INV_X4 u4_sub_472_U9 ( .A(u4_sub_472_carry_8_), .ZN(u4_sub_472_n4) );
  INV_X4 u4_sub_472_U8 ( .A(n4353), .ZN(u4_sub_472_n3) );
  XNOR2_X2 u4_sub_472_U7 ( .A(n4353), .B(u4_sub_472_carry_8_), .ZN(
        u4_exp_fix_diva[8]) );
  NAND2_X2 u4_sub_472_U6 ( .A1(u4_sub_472_n3), .A2(u4_sub_472_n4), .ZN(
        u4_sub_472_carry_9_) );
  INV_X4 u4_sub_472_U5 ( .A(u4_sub_472_carry_7_), .ZN(u4_sub_472_n2) );
  INV_X4 u4_sub_472_U4 ( .A(n4281), .ZN(u4_sub_472_n1) );
  XNOR2_X2 u4_sub_472_U3 ( .A(n4281), .B(u4_sub_472_carry_7_), .ZN(
        u4_exp_fix_diva[7]) );
  NAND2_X2 u4_sub_472_U2 ( .A1(u4_sub_472_n1), .A2(u4_sub_472_n2), .ZN(
        u4_sub_472_carry_8_) );
  XNOR2_X2 u4_sub_472_U1 ( .A(n4656), .B(u4_sub_472_carry_10_), .ZN(
        u4_exp_fix_diva[10]) );
  FA_X1 u4_sub_472_U2_1 ( .A(exp_r[1]), .B(u4_sub_472_n13), .CI(
        u4_sub_472_carry_1_), .CO(u4_sub_472_carry_2_), .S(u4_exp_fix_diva[1])
         );
  FA_X1 u4_sub_472_U2_2 ( .A(n4315), .B(u4_sub_472_n12), .CI(
        u4_sub_472_carry_2_), .CO(u4_sub_472_carry_3_), .S(u4_exp_fix_diva[2])
         );
  FA_X1 u4_sub_472_U2_3 ( .A(n4655), .B(u4_sub_472_n11), .CI(
        u4_sub_472_carry_3_), .CO(u4_sub_472_carry_4_), .S(u4_exp_fix_diva[3])
         );
  FA_X1 u4_sub_472_U2_4 ( .A(n4282), .B(u4_sub_472_n10), .CI(
        u4_sub_472_carry_4_), .CO(u4_sub_472_carry_5_), .S(u4_exp_fix_diva[4])
         );
  FA_X1 u4_sub_472_U2_5 ( .A(n4290), .B(u4_sub_472_n9), .CI(
        u4_sub_472_carry_5_), .CO(u4_sub_472_carry_6_), .S(u4_exp_fix_diva[5])
         );
  FA_X1 u4_sub_472_U2_6 ( .A(exp_r[6]), .B(u4_sub_472_n8), .CI(
        u4_sub_472_carry_6_), .CO(u4_sub_472_carry_7_), .S(u4_exp_fix_diva[6])
         );
  INV_X1 u4_add_464_U2 ( .A(u4_exp_out_0_), .ZN(u4_exp_out_pl1_0_) );
  XOR2_X1 u4_add_464_U1 ( .A(u4_add_464_carry[10]), .B(u4_exp_out_10_), .Z(
        u4_exp_out_pl1_10_) );
  HA_X1 u4_add_464_U1_1_1 ( .A(u4_exp_out_1_), .B(u4_exp_out_0_), .CO(
        u4_add_464_carry[2]), .S(u4_exp_out_pl1_1_) );
  HA_X1 u4_add_464_U1_1_2 ( .A(u4_exp_out_2_), .B(u4_add_464_carry[2]), .CO(
        u4_add_464_carry[3]), .S(u4_exp_out_pl1_2_) );
  HA_X1 u4_add_464_U1_1_3 ( .A(u4_exp_out_3_), .B(u4_add_464_carry[3]), .CO(
        u4_add_464_carry[4]), .S(u4_exp_out_pl1_3_) );
  HA_X1 u4_add_464_U1_1_4 ( .A(u4_exp_out_4_), .B(u4_add_464_carry[4]), .CO(
        u4_add_464_carry[5]), .S(u4_exp_out_pl1_4_) );
  HA_X1 u4_add_464_U1_1_5 ( .A(u4_exp_out_5_), .B(u4_add_464_carry[5]), .CO(
        u4_add_464_carry[6]), .S(u4_exp_out_pl1_5_) );
  HA_X1 u4_add_464_U1_1_6 ( .A(u4_exp_out_6_), .B(u4_add_464_carry[6]), .CO(
        u4_add_464_carry[7]), .S(u4_exp_out_pl1_6_) );
  HA_X1 u4_add_464_U1_1_7 ( .A(u4_exp_out_7_), .B(u4_add_464_carry[7]), .CO(
        u4_add_464_carry[8]), .S(u4_exp_out_pl1_7_) );
  HA_X1 u4_add_464_U1_1_8 ( .A(u4_exp_out_8_), .B(u4_add_464_carry[8]), .CO(
        u4_add_464_carry[9]), .S(u4_exp_out_pl1_8_) );
  HA_X1 u4_add_464_U1_1_9 ( .A(u4_exp_out_9_), .B(u4_add_464_carry[9]), .CO(
        u4_add_464_carry[10]), .S(u4_exp_out_pl1_9_) );
  INV_X1 u4_sll_454_U266 ( .A(u4_shift_left[8]), .ZN(u4_sll_454_n53) );
  OR2_X1 u4_sll_454_U265 ( .A1(u4_sll_454_n2), .A2(u4_shift_left[7]), .ZN(
        u4_sll_454_n85) );
  NAND2_X1 u4_sll_454_U264 ( .A1(u4_shift_left[7]), .A2(u4_sll_454_n3), .ZN(
        u4_sll_454_n87) );
  INV_X1 u4_sll_454_U263 ( .A(u4_sll_454_n87), .ZN(u4_sll_454_n86) );
  AOI21_X1 u4_sll_454_U262 ( .B1(u4_shift_left[0]), .B2(u4_sll_454_n85), .A(
        u4_sll_454_n86), .ZN(u4_sll_454_SHMAG_0_) );
  AND2_X1 u4_sll_454_U261 ( .A1(n6446), .A2(u4_sll_454_SHMAG_0_), .ZN(
        u4_sll_454_ML_int_1__0_) );
  AOI21_X1 u4_sll_454_U260 ( .B1(u4_shift_left[1]), .B2(u4_sll_454_n85), .A(
        u4_sll_454_n86), .ZN(u4_sll_454_SHMAG_1_) );
  AND2_X1 u4_sll_454_U259 ( .A1(u4_sll_454_ML_int_1__0_), .A2(
        u4_sll_454_SHMAG_1_), .ZN(u4_sll_454_ML_int_2__0_) );
  AND2_X1 u4_sll_454_U258 ( .A1(u4_sll_454_ML_int_1__1_), .A2(
        u4_sll_454_SHMAG_1_), .ZN(u4_sll_454_ML_int_2__1_) );
  AOI21_X1 u4_sll_454_U257 ( .B1(u4_shift_left[2]), .B2(u4_sll_454_n85), .A(
        u4_sll_454_n86), .ZN(u4_sll_454_SHMAG_2_) );
  AND2_X1 u4_sll_454_U256 ( .A1(u4_sll_454_ML_int_2__0_), .A2(
        u4_sll_454_SHMAG_2_), .ZN(u4_sll_454_ML_int_3__0_) );
  AND2_X1 u4_sll_454_U255 ( .A1(u4_sll_454_ML_int_2__1_), .A2(
        u4_sll_454_SHMAG_2_), .ZN(u4_sll_454_ML_int_3__1_) );
  AND2_X1 u4_sll_454_U254 ( .A1(u4_sll_454_ML_int_2__2_), .A2(
        u4_sll_454_SHMAG_2_), .ZN(u4_sll_454_ML_int_3__2_) );
  AND2_X1 u4_sll_454_U253 ( .A1(u4_sll_454_ML_int_2__3_), .A2(
        u4_sll_454_SHMAG_2_), .ZN(u4_sll_454_ML_int_3__3_) );
  AOI21_X1 u4_sll_454_U252 ( .B1(u4_shift_left[3]), .B2(u4_sll_454_n85), .A(
        u4_sll_454_n86), .ZN(u4_sll_454_SHMAG_3_) );
  AND2_X1 u4_sll_454_U251 ( .A1(u4_sll_454_ML_int_3__0_), .A2(u4_sll_454_n23), 
        .ZN(u4_sll_454_ML_int_4__0_) );
  AND2_X1 u4_sll_454_U250 ( .A1(u4_sll_454_ML_int_3__1_), .A2(u4_sll_454_n23), 
        .ZN(u4_sll_454_ML_int_4__1_) );
  AND2_X1 u4_sll_454_U249 ( .A1(u4_sll_454_ML_int_3__2_), .A2(u4_sll_454_n23), 
        .ZN(u4_sll_454_ML_int_4__2_) );
  AND2_X1 u4_sll_454_U248 ( .A1(u4_sll_454_ML_int_3__3_), .A2(u4_sll_454_n23), 
        .ZN(u4_sll_454_ML_int_4__3_) );
  AND2_X1 u4_sll_454_U247 ( .A1(u4_sll_454_ML_int_3__4_), .A2(u4_sll_454_n23), 
        .ZN(u4_sll_454_ML_int_4__4_) );
  AND2_X1 u4_sll_454_U246 ( .A1(u4_sll_454_ML_int_3__5_), .A2(u4_sll_454_n23), 
        .ZN(u4_sll_454_ML_int_4__5_) );
  AND2_X1 u4_sll_454_U245 ( .A1(u4_sll_454_ML_int_3__6_), .A2(u4_sll_454_n23), 
        .ZN(u4_sll_454_ML_int_4__6_) );
  AND2_X1 u4_sll_454_U244 ( .A1(u4_sll_454_ML_int_3__7_), .A2(u4_sll_454_n23), 
        .ZN(u4_sll_454_ML_int_4__7_) );
  AOI21_X1 u4_sll_454_U243 ( .B1(u4_shift_left[4]), .B2(u4_sll_454_n85), .A(
        u4_sll_454_n86), .ZN(u4_sll_454_SHMAG_4_) );
  AND2_X1 u4_sll_454_U242 ( .A1(u4_sll_454_ML_int_4__0_), .A2(u4_sll_454_n35), 
        .ZN(u4_sll_454_ML_int_5__0_) );
  AND2_X1 u4_sll_454_U241 ( .A1(u4_sll_454_ML_int_4__10_), .A2(u4_sll_454_n25), 
        .ZN(u4_sll_454_ML_int_5__10_) );
  AND2_X1 u4_sll_454_U240 ( .A1(u4_sll_454_ML_int_4__11_), .A2(u4_sll_454_n25), 
        .ZN(u4_sll_454_ML_int_5__11_) );
  AND2_X1 u4_sll_454_U239 ( .A1(u4_sll_454_ML_int_4__12_), .A2(u4_sll_454_n25), 
        .ZN(u4_sll_454_ML_int_5__12_) );
  AND2_X1 u4_sll_454_U238 ( .A1(u4_sll_454_ML_int_4__13_), .A2(u4_sll_454_n25), 
        .ZN(u4_sll_454_ML_int_5__13_) );
  AND2_X1 u4_sll_454_U237 ( .A1(u4_sll_454_ML_int_4__14_), .A2(u4_sll_454_n25), 
        .ZN(u4_sll_454_ML_int_5__14_) );
  AND2_X1 u4_sll_454_U236 ( .A1(u4_sll_454_ML_int_4__15_), .A2(u4_sll_454_n25), 
        .ZN(u4_sll_454_ML_int_5__15_) );
  AND2_X1 u4_sll_454_U235 ( .A1(u4_sll_454_ML_int_4__1_), .A2(u4_sll_454_n35), 
        .ZN(u4_sll_454_ML_int_5__1_) );
  AND2_X1 u4_sll_454_U234 ( .A1(u4_sll_454_ML_int_4__2_), .A2(u4_sll_454_n26), 
        .ZN(u4_sll_454_ML_int_5__2_) );
  AND2_X1 u4_sll_454_U233 ( .A1(u4_sll_454_ML_int_4__3_), .A2(u4_sll_454_n26), 
        .ZN(u4_sll_454_ML_int_5__3_) );
  AND2_X1 u4_sll_454_U232 ( .A1(u4_sll_454_ML_int_4__4_), .A2(u4_sll_454_n26), 
        .ZN(u4_sll_454_ML_int_5__4_) );
  AND2_X1 u4_sll_454_U231 ( .A1(u4_sll_454_ML_int_4__5_), .A2(u4_sll_454_n26), 
        .ZN(u4_sll_454_ML_int_5__5_) );
  AND2_X1 u4_sll_454_U230 ( .A1(u4_sll_454_ML_int_4__6_), .A2(u4_sll_454_n26), 
        .ZN(u4_sll_454_ML_int_5__6_) );
  AND2_X1 u4_sll_454_U229 ( .A1(u4_sll_454_ML_int_4__7_), .A2(u4_sll_454_n26), 
        .ZN(u4_sll_454_ML_int_5__7_) );
  AND2_X1 u4_sll_454_U228 ( .A1(u4_sll_454_ML_int_4__8_), .A2(u4_sll_454_n26), 
        .ZN(u4_sll_454_ML_int_5__8_) );
  AND2_X1 u4_sll_454_U227 ( .A1(u4_sll_454_ML_int_4__9_), .A2(u4_sll_454_n26), 
        .ZN(u4_sll_454_ML_int_5__9_) );
  NAND2_X1 u4_sll_454_U226 ( .A1(u4_shift_left[5]), .A2(u4_sll_454_n85), .ZN(
        u4_sll_454_n88) );
  NAND2_X1 u4_sll_454_U225 ( .A1(u4_sll_454_n87), .A2(u4_sll_454_n88), .ZN(
        u4_sll_454_temp_int_SH_5_) );
  NAND2_X1 u4_sll_454_U224 ( .A1(u4_sll_454_ML_int_5__0_), .A2(u4_sll_454_n39), 
        .ZN(u4_sll_454_n84) );
  INV_X1 u4_sll_454_U223 ( .A(u4_sll_454_n84), .ZN(u4_sll_454_ML_int_6__0_) );
  NAND2_X1 u4_sll_454_U222 ( .A1(u4_sll_454_ML_int_5__10_), .A2(u4_sll_454_n39), .ZN(u4_sll_454_n83) );
  INV_X1 u4_sll_454_U221 ( .A(u4_sll_454_n83), .ZN(u4_sll_454_ML_int_6__10_)
         );
  NAND2_X1 u4_sll_454_U220 ( .A1(u4_sll_454_ML_int_5__11_), .A2(u4_sll_454_n39), .ZN(u4_sll_454_n82) );
  INV_X1 u4_sll_454_U219 ( .A(u4_sll_454_n82), .ZN(u4_sll_454_ML_int_6__11_)
         );
  NAND2_X1 u4_sll_454_U218 ( .A1(u4_sll_454_ML_int_5__12_), .A2(u4_sll_454_n40), .ZN(u4_sll_454_n81) );
  INV_X1 u4_sll_454_U217 ( .A(u4_sll_454_n81), .ZN(u4_sll_454_ML_int_6__12_)
         );
  NAND2_X1 u4_sll_454_U216 ( .A1(u4_sll_454_ML_int_5__13_), .A2(u4_sll_454_n39), .ZN(u4_sll_454_n80) );
  INV_X1 u4_sll_454_U215 ( .A(u4_sll_454_n80), .ZN(u4_sll_454_ML_int_6__13_)
         );
  NAND2_X1 u4_sll_454_U214 ( .A1(u4_sll_454_ML_int_5__14_), .A2(u4_sll_454_n40), .ZN(u4_sll_454_n79) );
  INV_X1 u4_sll_454_U213 ( .A(u4_sll_454_n79), .ZN(u4_sll_454_ML_int_6__14_)
         );
  NAND2_X1 u4_sll_454_U212 ( .A1(u4_sll_454_ML_int_5__15_), .A2(u4_sll_454_n40), .ZN(u4_sll_454_n78) );
  INV_X1 u4_sll_454_U211 ( .A(u4_sll_454_n78), .ZN(u4_sll_454_ML_int_6__15_)
         );
  NAND2_X1 u4_sll_454_U210 ( .A1(u4_sll_454_ML_int_5__16_), .A2(u4_sll_454_n40), .ZN(u4_sll_454_n77) );
  INV_X1 u4_sll_454_U209 ( .A(u4_sll_454_n77), .ZN(u4_sll_454_ML_int_6__16_)
         );
  NAND2_X1 u4_sll_454_U208 ( .A1(u4_sll_454_ML_int_5__17_), .A2(u4_sll_454_n40), .ZN(u4_sll_454_n76) );
  INV_X1 u4_sll_454_U207 ( .A(u4_sll_454_n76), .ZN(u4_sll_454_ML_int_6__17_)
         );
  NAND2_X1 u4_sll_454_U206 ( .A1(u4_sll_454_ML_int_5__18_), .A2(u4_sll_454_n40), .ZN(u4_sll_454_n75) );
  INV_X1 u4_sll_454_U205 ( .A(u4_sll_454_n75), .ZN(u4_sll_454_ML_int_6__18_)
         );
  NAND2_X1 u4_sll_454_U204 ( .A1(u4_sll_454_ML_int_5__19_), .A2(u4_sll_454_n40), .ZN(u4_sll_454_n74) );
  INV_X1 u4_sll_454_U203 ( .A(u4_sll_454_n74), .ZN(u4_sll_454_ML_int_6__19_)
         );
  NAND2_X1 u4_sll_454_U202 ( .A1(u4_sll_454_ML_int_5__1_), .A2(u4_sll_454_n41), 
        .ZN(u4_sll_454_n73) );
  INV_X1 u4_sll_454_U201 ( .A(u4_sll_454_n73), .ZN(u4_sll_454_ML_int_6__1_) );
  NAND2_X1 u4_sll_454_U200 ( .A1(u4_sll_454_ML_int_5__20_), .A2(u4_sll_454_n40), .ZN(u4_sll_454_n72) );
  INV_X1 u4_sll_454_U199 ( .A(u4_sll_454_n72), .ZN(u4_sll_454_ML_int_6__20_)
         );
  NAND2_X1 u4_sll_454_U198 ( .A1(u4_sll_454_ML_int_5__21_), .A2(u4_sll_454_n40), .ZN(u4_sll_454_n71) );
  INV_X1 u4_sll_454_U197 ( .A(u4_sll_454_n71), .ZN(u4_sll_454_ML_int_6__21_)
         );
  NAND2_X1 u4_sll_454_U196 ( .A1(u4_sll_454_ML_int_5__22_), .A2(u4_sll_454_n40), .ZN(u4_sll_454_n70) );
  INV_X1 u4_sll_454_U195 ( .A(u4_sll_454_n70), .ZN(u4_sll_454_ML_int_6__22_)
         );
  NAND2_X1 u4_sll_454_U194 ( .A1(u4_sll_454_ML_int_5__23_), .A2(u4_sll_454_n40), .ZN(u4_sll_454_n69) );
  INV_X1 u4_sll_454_U193 ( .A(u4_sll_454_n69), .ZN(u4_sll_454_ML_int_6__23_)
         );
  NAND2_X1 u4_sll_454_U192 ( .A1(u4_sll_454_ML_int_5__24_), .A2(u4_sll_454_n40), .ZN(u4_sll_454_n68) );
  INV_X1 u4_sll_454_U191 ( .A(u4_sll_454_n68), .ZN(u4_sll_454_ML_int_6__24_)
         );
  NAND2_X1 u4_sll_454_U190 ( .A1(u4_sll_454_ML_int_5__25_), .A2(u4_sll_454_n40), .ZN(u4_sll_454_n67) );
  INV_X1 u4_sll_454_U189 ( .A(u4_sll_454_n67), .ZN(u4_sll_454_ML_int_6__25_)
         );
  NAND2_X1 u4_sll_454_U188 ( .A1(u4_sll_454_ML_int_5__26_), .A2(u4_sll_454_n41), .ZN(u4_sll_454_n66) );
  INV_X1 u4_sll_454_U187 ( .A(u4_sll_454_n66), .ZN(u4_sll_454_ML_int_6__26_)
         );
  NAND2_X1 u4_sll_454_U186 ( .A1(u4_sll_454_ML_int_5__27_), .A2(u4_sll_454_n41), .ZN(u4_sll_454_n65) );
  INV_X1 u4_sll_454_U185 ( .A(u4_sll_454_n65), .ZN(u4_sll_454_ML_int_6__27_)
         );
  NAND2_X1 u4_sll_454_U184 ( .A1(u4_sll_454_ML_int_5__28_), .A2(u4_sll_454_n41), .ZN(u4_sll_454_n64) );
  INV_X1 u4_sll_454_U183 ( .A(u4_sll_454_n64), .ZN(u4_sll_454_ML_int_6__28_)
         );
  NAND2_X1 u4_sll_454_U182 ( .A1(u4_sll_454_ML_int_5__29_), .A2(u4_sll_454_n41), .ZN(u4_sll_454_n63) );
  INV_X1 u4_sll_454_U181 ( .A(u4_sll_454_n63), .ZN(u4_sll_454_ML_int_6__29_)
         );
  NAND2_X1 u4_sll_454_U180 ( .A1(u4_sll_454_ML_int_5__2_), .A2(u4_sll_454_n41), 
        .ZN(u4_sll_454_n62) );
  INV_X1 u4_sll_454_U179 ( .A(u4_sll_454_n62), .ZN(u4_sll_454_ML_int_6__2_) );
  NAND2_X1 u4_sll_454_U178 ( .A1(u4_sll_454_ML_int_5__30_), .A2(u4_sll_454_n41), .ZN(u4_sll_454_n61) );
  INV_X1 u4_sll_454_U177 ( .A(u4_sll_454_n61), .ZN(u4_sll_454_ML_int_6__30_)
         );
  NAND2_X1 u4_sll_454_U176 ( .A1(u4_sll_454_ML_int_5__31_), .A2(u4_sll_454_n41), .ZN(u4_sll_454_n60) );
  INV_X1 u4_sll_454_U175 ( .A(u4_sll_454_n60), .ZN(u4_sll_454_ML_int_6__31_)
         );
  NAND2_X1 u4_sll_454_U174 ( .A1(u4_sll_454_ML_int_5__3_), .A2(u4_sll_454_n41), 
        .ZN(u4_sll_454_n59) );
  INV_X1 u4_sll_454_U173 ( .A(u4_sll_454_n59), .ZN(u4_sll_454_ML_int_6__3_) );
  NAND2_X1 u4_sll_454_U172 ( .A1(u4_sll_454_ML_int_5__4_), .A2(u4_sll_454_n41), 
        .ZN(u4_sll_454_n58) );
  INV_X1 u4_sll_454_U171 ( .A(u4_sll_454_n58), .ZN(u4_sll_454_ML_int_6__4_) );
  NAND2_X1 u4_sll_454_U170 ( .A1(u4_sll_454_ML_int_5__5_), .A2(u4_sll_454_n41), 
        .ZN(u4_sll_454_n57) );
  INV_X1 u4_sll_454_U169 ( .A(u4_sll_454_n57), .ZN(u4_sll_454_ML_int_6__5_) );
  NAND2_X1 u4_sll_454_U168 ( .A1(u4_sll_454_ML_int_5__6_), .A2(u4_sll_454_n41), 
        .ZN(u4_sll_454_n56) );
  INV_X1 u4_sll_454_U167 ( .A(u4_sll_454_n56), .ZN(u4_sll_454_ML_int_6__6_) );
  NAND2_X1 u4_sll_454_U166 ( .A1(u4_sll_454_ML_int_5__7_), .A2(u4_sll_454_n41), 
        .ZN(u4_sll_454_n55) );
  INV_X1 u4_sll_454_U165 ( .A(u4_sll_454_n55), .ZN(u4_sll_454_ML_int_6__7_) );
  NAND2_X1 u4_sll_454_U164 ( .A1(u4_sll_454_ML_int_5__8_), .A2(u4_sll_454_n41), 
        .ZN(u4_sll_454_n54) );
  INV_X1 u4_sll_454_U163 ( .A(u4_sll_454_n54), .ZN(u4_sll_454_ML_int_6__8_) );
  NAND2_X1 u4_sll_454_U162 ( .A1(u4_sll_454_ML_int_5__9_), .A2(u4_sll_454_n41), 
        .ZN(u4_sll_454_n52) );
  INV_X1 u4_sll_454_U161 ( .A(u4_sll_454_n52), .ZN(u4_sll_454_ML_int_6__9_) );
  AOI21_X1 u4_sll_454_U160 ( .B1(u4_shift_left[6]), .B2(u4_sll_454_n85), .A(
        u4_sll_454_n86), .ZN(u4_sll_454_SHMAG_6_) );
  NOR2_X1 u4_sll_454_U159 ( .A1(u4_sll_454_n4), .A2(u4_sll_454_n84), .ZN(
        u4_N6014) );
  AND2_X1 u4_sll_454_U158 ( .A1(u4_sll_454_ML_int_7__100_), .A2(u4_sll_454_n3), 
        .ZN(u4_N6114) );
  AND2_X1 u4_sll_454_U157 ( .A1(u4_sll_454_ML_int_7__101_), .A2(u4_sll_454_n3), 
        .ZN(u4_N6115) );
  AND2_X1 u4_sll_454_U156 ( .A1(u4_sll_454_ML_int_7__102_), .A2(u4_sll_454_n3), 
        .ZN(u4_N6116) );
  AND2_X1 u4_sll_454_U155 ( .A1(u4_sll_454_ML_int_7__103_), .A2(u4_sll_454_n3), 
        .ZN(u4_N6117) );
  AND2_X1 u4_sll_454_U154 ( .A1(u4_sll_454_ML_int_7__104_), .A2(u4_sll_454_n3), 
        .ZN(u4_N6118) );
  AND2_X1 u4_sll_454_U153 ( .A1(u4_sll_454_ML_int_7__105_), .A2(u4_sll_454_n3), 
        .ZN(u4_N6119) );
  NOR2_X1 u4_sll_454_U152 ( .A1(u4_sll_454_n4), .A2(u4_sll_454_n83), .ZN(
        u4_N6024) );
  NOR2_X1 u4_sll_454_U151 ( .A1(u4_sll_454_n4), .A2(u4_sll_454_n82), .ZN(
        u4_N6025) );
  NOR2_X1 u4_sll_454_U150 ( .A1(u4_sll_454_n4), .A2(u4_sll_454_n81), .ZN(
        u4_N6026) );
  NOR2_X1 u4_sll_454_U149 ( .A1(u4_sll_454_n4), .A2(u4_sll_454_n80), .ZN(
        u4_N6027) );
  NOR2_X1 u4_sll_454_U148 ( .A1(u4_sll_454_n4), .A2(u4_sll_454_n79), .ZN(
        u4_N6028) );
  NOR2_X1 u4_sll_454_U147 ( .A1(u4_sll_454_n4), .A2(u4_sll_454_n78), .ZN(
        u4_N6029) );
  NOR2_X1 u4_sll_454_U146 ( .A1(u4_sll_454_n4), .A2(u4_sll_454_n77), .ZN(
        u4_N6030) );
  NOR2_X1 u4_sll_454_U145 ( .A1(u4_sll_454_n4), .A2(u4_sll_454_n76), .ZN(
        u4_N6031) );
  NOR2_X1 u4_sll_454_U144 ( .A1(u4_sll_454_n4), .A2(u4_sll_454_n75), .ZN(
        u4_N6032) );
  NOR2_X1 u4_sll_454_U143 ( .A1(u4_sll_454_n4), .A2(u4_sll_454_n74), .ZN(
        u4_N6033) );
  NOR2_X1 u4_sll_454_U142 ( .A1(u4_sll_454_n5), .A2(u4_sll_454_n73), .ZN(
        u4_N6015) );
  NOR2_X1 u4_sll_454_U141 ( .A1(u4_sll_454_n5), .A2(u4_sll_454_n72), .ZN(
        u4_N6034) );
  NOR2_X1 u4_sll_454_U140 ( .A1(u4_sll_454_n5), .A2(u4_sll_454_n71), .ZN(
        u4_N6035) );
  NOR2_X1 u4_sll_454_U139 ( .A1(u4_sll_454_n5), .A2(u4_sll_454_n70), .ZN(
        u4_N6036) );
  NOR2_X1 u4_sll_454_U138 ( .A1(u4_sll_454_n5), .A2(u4_sll_454_n69), .ZN(
        u4_N6037) );
  NOR2_X1 u4_sll_454_U137 ( .A1(u4_sll_454_n5), .A2(u4_sll_454_n68), .ZN(
        u4_N6038) );
  NOR2_X1 u4_sll_454_U136 ( .A1(u4_sll_454_n5), .A2(u4_sll_454_n67), .ZN(
        u4_N6039) );
  NOR2_X1 u4_sll_454_U135 ( .A1(u4_sll_454_n5), .A2(u4_sll_454_n66), .ZN(
        u4_N6040) );
  NOR2_X1 u4_sll_454_U134 ( .A1(u4_sll_454_n5), .A2(u4_sll_454_n65), .ZN(
        u4_N6041) );
  NOR2_X1 u4_sll_454_U133 ( .A1(u4_sll_454_n5), .A2(u4_sll_454_n64), .ZN(
        u4_N6042) );
  NOR2_X1 u4_sll_454_U132 ( .A1(u4_sll_454_n5), .A2(u4_sll_454_n63), .ZN(
        u4_N6043) );
  NOR2_X1 u4_sll_454_U131 ( .A1(u4_sll_454_n4), .A2(u4_sll_454_n62), .ZN(
        u4_N6016) );
  NOR2_X1 u4_sll_454_U130 ( .A1(u4_sll_454_n4), .A2(u4_sll_454_n61), .ZN(
        u4_N6044) );
  NOR2_X1 u4_sll_454_U129 ( .A1(u4_sll_454_n5), .A2(u4_sll_454_n60), .ZN(
        u4_N6045) );
  AND2_X1 u4_sll_454_U128 ( .A1(u4_sll_454_ML_int_6__32_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6046) );
  AND2_X1 u4_sll_454_U127 ( .A1(u4_sll_454_ML_int_6__33_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6047) );
  AND2_X1 u4_sll_454_U126 ( .A1(u4_sll_454_ML_int_6__34_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6048) );
  AND2_X1 u4_sll_454_U125 ( .A1(u4_sll_454_ML_int_6__35_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6049) );
  AND2_X1 u4_sll_454_U124 ( .A1(u4_sll_454_ML_int_6__36_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6050) );
  AND2_X1 u4_sll_454_U123 ( .A1(u4_sll_454_ML_int_6__37_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6051) );
  AND2_X1 u4_sll_454_U122 ( .A1(u4_sll_454_ML_int_6__38_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6052) );
  AND2_X1 u4_sll_454_U121 ( .A1(u4_sll_454_ML_int_6__39_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6053) );
  NOR2_X1 u4_sll_454_U120 ( .A1(u4_sll_454_n4), .A2(u4_sll_454_n59), .ZN(
        u4_N6017) );
  AND2_X1 u4_sll_454_U119 ( .A1(u4_sll_454_ML_int_6__40_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6054) );
  AND2_X1 u4_sll_454_U118 ( .A1(u4_sll_454_ML_int_6__41_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6055) );
  AND2_X1 u4_sll_454_U117 ( .A1(u4_sll_454_ML_int_6__42_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6056) );
  AND2_X1 u4_sll_454_U116 ( .A1(u4_sll_454_ML_int_6__43_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6057) );
  AND2_X1 u4_sll_454_U115 ( .A1(u4_sll_454_ML_int_6__44_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6058) );
  AND2_X1 u4_sll_454_U114 ( .A1(u4_sll_454_ML_int_6__45_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6059) );
  AND2_X1 u4_sll_454_U113 ( .A1(u4_sll_454_ML_int_6__46_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6060) );
  AND2_X1 u4_sll_454_U112 ( .A1(u4_sll_454_ML_int_6__47_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6061) );
  AND2_X1 u4_sll_454_U111 ( .A1(u4_sll_454_ML_int_6__48_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6062) );
  AND2_X1 u4_sll_454_U110 ( .A1(u4_sll_454_ML_int_6__49_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6063) );
  NOR2_X1 u4_sll_454_U109 ( .A1(u4_sll_454_n4), .A2(u4_sll_454_n58), .ZN(
        u4_N6018) );
  AND2_X1 u4_sll_454_U108 ( .A1(u4_sll_454_ML_int_6__50_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6064) );
  AND2_X1 u4_sll_454_U107 ( .A1(u4_sll_454_ML_int_6__51_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6065) );
  AND2_X1 u4_sll_454_U106 ( .A1(u4_sll_454_ML_int_6__52_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6066) );
  AND2_X1 u4_sll_454_U105 ( .A1(u4_sll_454_ML_int_6__53_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6067) );
  AND2_X1 u4_sll_454_U104 ( .A1(u4_sll_454_ML_int_6__54_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6068) );
  AND2_X1 u4_sll_454_U103 ( .A1(u4_sll_454_ML_int_6__55_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6069) );
  AND2_X1 u4_sll_454_U102 ( .A1(u4_sll_454_ML_int_6__56_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6070) );
  AND2_X1 u4_sll_454_U101 ( .A1(u4_sll_454_ML_int_6__57_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6071) );
  AND2_X1 u4_sll_454_U100 ( .A1(u4_sll_454_ML_int_6__58_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6072) );
  AND2_X1 u4_sll_454_U99 ( .A1(u4_sll_454_ML_int_6__59_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6073) );
  NOR2_X1 u4_sll_454_U98 ( .A1(u4_sll_454_n4), .A2(u4_sll_454_n57), .ZN(
        u4_N6019) );
  AND2_X1 u4_sll_454_U97 ( .A1(u4_sll_454_ML_int_6__60_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6074) );
  AND2_X1 u4_sll_454_U96 ( .A1(u4_sll_454_ML_int_6__61_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6075) );
  AND2_X1 u4_sll_454_U95 ( .A1(u4_sll_454_ML_int_6__62_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6076) );
  AND2_X1 u4_sll_454_U94 ( .A1(u4_sll_454_ML_int_6__63_), .A2(u4_sll_454_n1), 
        .ZN(u4_N6077) );
  AND2_X1 u4_sll_454_U93 ( .A1(u4_sll_454_ML_int_7__64_), .A2(u4_sll_454_n3), 
        .ZN(u4_N6078) );
  AND2_X1 u4_sll_454_U92 ( .A1(u4_sll_454_ML_int_7__65_), .A2(u4_sll_454_n3), 
        .ZN(u4_N6079) );
  AND2_X1 u4_sll_454_U91 ( .A1(u4_sll_454_ML_int_7__66_), .A2(u4_sll_454_n3), 
        .ZN(u4_N6080) );
  AND2_X1 u4_sll_454_U90 ( .A1(u4_sll_454_ML_int_7__67_), .A2(u4_sll_454_n3), 
        .ZN(u4_N6081) );
  AND2_X1 u4_sll_454_U89 ( .A1(u4_sll_454_ML_int_7__68_), .A2(u4_sll_454_n2), 
        .ZN(u4_N6082) );
  AND2_X1 u4_sll_454_U88 ( .A1(u4_sll_454_ML_int_7__69_), .A2(u4_sll_454_n2), 
        .ZN(u4_N6083) );
  NOR2_X1 u4_sll_454_U87 ( .A1(u4_sll_454_n4), .A2(u4_sll_454_n56), .ZN(
        u4_N6020) );
  AND2_X1 u4_sll_454_U86 ( .A1(u4_sll_454_ML_int_7__70_), .A2(u4_sll_454_n53), 
        .ZN(u4_N6084) );
  AND2_X1 u4_sll_454_U85 ( .A1(u4_sll_454_ML_int_7__71_), .A2(u4_sll_454_n53), 
        .ZN(u4_N6085) );
  AND2_X1 u4_sll_454_U84 ( .A1(u4_sll_454_ML_int_7__72_), .A2(u4_sll_454_n53), 
        .ZN(u4_N6086) );
  AND2_X1 u4_sll_454_U83 ( .A1(u4_sll_454_ML_int_7__73_), .A2(u4_sll_454_n53), 
        .ZN(u4_N6087) );
  AND2_X1 u4_sll_454_U82 ( .A1(u4_sll_454_ML_int_7__74_), .A2(u4_sll_454_n53), 
        .ZN(u4_N6088) );
  AND2_X1 u4_sll_454_U81 ( .A1(u4_sll_454_ML_int_7__75_), .A2(u4_sll_454_n53), 
        .ZN(u4_N6089) );
  AND2_X1 u4_sll_454_U80 ( .A1(u4_sll_454_ML_int_7__76_), .A2(u4_sll_454_n53), 
        .ZN(u4_N6090) );
  AND2_X1 u4_sll_454_U79 ( .A1(u4_sll_454_ML_int_7__77_), .A2(u4_sll_454_n53), 
        .ZN(u4_N6091) );
  AND2_X1 u4_sll_454_U78 ( .A1(u4_sll_454_ML_int_7__78_), .A2(u4_sll_454_n53), 
        .ZN(u4_N6092) );
  AND2_X1 u4_sll_454_U77 ( .A1(u4_sll_454_ML_int_7__79_), .A2(u4_sll_454_n53), 
        .ZN(u4_N6093) );
  NOR2_X1 u4_sll_454_U76 ( .A1(u4_sll_454_n5), .A2(u4_sll_454_n55), .ZN(
        u4_N6021) );
  AND2_X1 u4_sll_454_U75 ( .A1(u4_sll_454_ML_int_7__80_), .A2(u4_sll_454_n53), 
        .ZN(u4_N6094) );
  AND2_X1 u4_sll_454_U74 ( .A1(u4_sll_454_ML_int_7__81_), .A2(u4_sll_454_n53), 
        .ZN(u4_N6095) );
  AND2_X1 u4_sll_454_U73 ( .A1(u4_sll_454_ML_int_7__82_), .A2(u4_sll_454_n53), 
        .ZN(u4_N6096) );
  AND2_X1 u4_sll_454_U72 ( .A1(u4_sll_454_ML_int_7__83_), .A2(u4_sll_454_n53), 
        .ZN(u4_N6097) );
  AND2_X1 u4_sll_454_U71 ( .A1(u4_sll_454_ML_int_7__84_), .A2(u4_sll_454_n53), 
        .ZN(u4_N6098) );
  AND2_X1 u4_sll_454_U70 ( .A1(u4_sll_454_ML_int_7__85_), .A2(u4_sll_454_n53), 
        .ZN(u4_N6099) );
  AND2_X1 u4_sll_454_U69 ( .A1(u4_sll_454_ML_int_7__86_), .A2(u4_sll_454_n53), 
        .ZN(u4_N6100) );
  AND2_X1 u4_sll_454_U68 ( .A1(u4_sll_454_ML_int_7__87_), .A2(u4_sll_454_n53), 
        .ZN(u4_N6101) );
  AND2_X1 u4_sll_454_U67 ( .A1(u4_sll_454_ML_int_7__88_), .A2(u4_sll_454_n53), 
        .ZN(u4_N6102) );
  AND2_X1 u4_sll_454_U66 ( .A1(u4_sll_454_ML_int_7__89_), .A2(u4_sll_454_n2), 
        .ZN(u4_N6103) );
  NOR2_X1 u4_sll_454_U65 ( .A1(u4_sll_454_n4), .A2(u4_sll_454_n54), .ZN(
        u4_N6022) );
  AND2_X1 u4_sll_454_U64 ( .A1(u4_sll_454_ML_int_7__90_), .A2(u4_sll_454_n2), 
        .ZN(u4_N6104) );
  AND2_X1 u4_sll_454_U63 ( .A1(u4_sll_454_ML_int_7__91_), .A2(u4_sll_454_n2), 
        .ZN(u4_N6105) );
  AND2_X1 u4_sll_454_U62 ( .A1(u4_sll_454_ML_int_7__92_), .A2(u4_sll_454_n2), 
        .ZN(u4_N6106) );
  AND2_X1 u4_sll_454_U61 ( .A1(u4_sll_454_ML_int_7__93_), .A2(u4_sll_454_n2), 
        .ZN(u4_N6107) );
  AND2_X1 u4_sll_454_U60 ( .A1(u4_sll_454_ML_int_7__94_), .A2(u4_sll_454_n2), 
        .ZN(u4_N6108) );
  AND2_X1 u4_sll_454_U59 ( .A1(u4_sll_454_ML_int_7__95_), .A2(u4_sll_454_n2), 
        .ZN(u4_N6109) );
  AND2_X1 u4_sll_454_U58 ( .A1(u4_sll_454_ML_int_7__96_), .A2(u4_sll_454_n2), 
        .ZN(u4_N6110) );
  AND2_X1 u4_sll_454_U57 ( .A1(u4_sll_454_ML_int_7__97_), .A2(u4_sll_454_n2), 
        .ZN(u4_N6111) );
  AND2_X1 u4_sll_454_U56 ( .A1(u4_sll_454_ML_int_7__98_), .A2(u4_sll_454_n2), 
        .ZN(u4_N6112) );
  AND2_X1 u4_sll_454_U55 ( .A1(u4_sll_454_ML_int_7__99_), .A2(u4_sll_454_n2), 
        .ZN(u4_N6113) );
  NOR2_X1 u4_sll_454_U54 ( .A1(u4_sll_454_n4), .A2(u4_sll_454_n52), .ZN(
        u4_N6023) );
  INV_X4 u4_sll_454_U53 ( .A(u4_sll_454_n1), .ZN(u4_sll_454_n5) );
  INV_X4 u4_sll_454_U52 ( .A(u4_sll_454_n1), .ZN(u4_sll_454_n4) );
  INV_X4 u4_sll_454_U51 ( .A(u4_sll_454_n39), .ZN(u4_sll_454_n43) );
  INV_X4 u4_sll_454_U50 ( .A(u4_sll_454_n50), .ZN(u4_sll_454_n48) );
  INV_X4 u4_sll_454_U49 ( .A(u4_sll_454_n35), .ZN(u4_sll_454_n28) );
  INV_X4 u4_sll_454_U48 ( .A(u4_sll_454_SHMAG_2_), .ZN(u4_sll_454_n15) );
  INV_X4 u4_sll_454_U47 ( .A(u4_sll_454_n39), .ZN(u4_sll_454_n42) );
  INV_X4 u4_sll_454_U46 ( .A(u4_sll_454_n35), .ZN(u4_sll_454_n27) );
  INV_X4 u4_sll_454_U45 ( .A(u4_sll_454_n24), .ZN(u4_sll_454_n23) );
  INV_X4 u4_sll_454_U44 ( .A(u4_sll_454_SHMAG_0_), .ZN(u4_sll_454_n8) );
  INV_X4 u4_sll_454_U43 ( .A(u4_sll_454_SHMAG_6_), .ZN(u4_sll_454_n38) );
  INV_X4 u4_sll_454_U42 ( .A(u4_sll_454_SHMAG_6_), .ZN(u4_sll_454_n37) );
  INV_X4 u4_sll_454_U41 ( .A(u4_sll_454_n27), .ZN(u4_sll_454_n25) );
  INV_X4 u4_sll_454_U40 ( .A(u4_sll_454_n23), .ZN(u4_sll_454_n18) );
  INV_X4 u4_sll_454_U39 ( .A(u4_sll_454_SHMAG_1_), .ZN(u4_sll_454_n11) );
  INV_X4 u4_sll_454_U38 ( .A(u4_sll_454_SHMAG_0_), .ZN(u4_sll_454_n7) );
  INV_X4 u4_sll_454_U37 ( .A(u4_shift_left[8]), .ZN(u4_sll_454_n3) );
  INV_X4 u4_sll_454_U36 ( .A(u4_shift_left[8]), .ZN(u4_sll_454_n2) );
  INV_X4 u4_sll_454_U35 ( .A(u4_sll_454_SHMAG_2_), .ZN(u4_sll_454_n14) );
  INV_X4 u4_sll_454_U34 ( .A(u4_sll_454_n36), .ZN(u4_sll_454_n35) );
  INV_X4 u4_sll_454_U33 ( .A(u4_sll_454_SHMAG_0_), .ZN(u4_sll_454_n6) );
  INV_X4 u4_sll_454_U32 ( .A(u4_sll_454_n47), .ZN(u4_sll_454_n39) );
  INV_X4 u4_sll_454_U31 ( .A(u4_sll_454_n49), .ZN(u4_sll_454_n44) );
  INV_X4 u4_sll_454_U30 ( .A(u4_sll_454_n36), .ZN(u4_sll_454_n33) );
  INV_X4 u4_sll_454_U29 ( .A(u4_sll_454_SHMAG_0_), .ZN(u4_sll_454_n9) );
  NOR2_X2 u4_sll_454_U28 ( .A1(u4_sll_454_n37), .A2(u4_shift_left[8]), .ZN(
        u4_sll_454_n1) );
  INV_X4 u4_sll_454_U27 ( .A(u4_sll_454_n43), .ZN(u4_sll_454_n40) );
  INV_X4 u4_sll_454_U26 ( .A(u4_sll_454_SHMAG_1_), .ZN(u4_sll_454_n10) );
  INV_X4 u4_sll_454_U25 ( .A(u4_sll_454_SHMAG_1_), .ZN(u4_sll_454_n13) );
  INV_X4 u4_sll_454_U24 ( .A(u4_sll_454_SHMAG_1_), .ZN(u4_sll_454_n12) );
  INV_X4 u4_sll_454_U23 ( .A(u4_sll_454_SHMAG_2_), .ZN(u4_sll_454_n17) );
  INV_X4 u4_sll_454_U22 ( .A(u4_sll_454_SHMAG_2_), .ZN(u4_sll_454_n16) );
  INV_X4 u4_sll_454_U21 ( .A(u4_sll_454_n36), .ZN(u4_sll_454_n34) );
  INV_X4 u4_sll_454_U20 ( .A(u4_sll_454_n51), .ZN(u4_sll_454_n50) );
  INV_X4 u4_sll_454_U19 ( .A(u4_sll_454_n48), .ZN(u4_sll_454_n47) );
  INV_X4 u4_sll_454_U18 ( .A(u4_sll_454_n50), .ZN(u4_sll_454_n49) );
  INV_X4 u4_sll_454_U17 ( .A(u4_sll_454_n28), .ZN(u4_sll_454_n26) );
  INV_X4 u4_sll_454_U16 ( .A(u4_sll_454_n42), .ZN(u4_sll_454_n41) );
  INV_X4 u4_sll_454_U15 ( .A(u4_sll_454_n23), .ZN(u4_sll_454_n19) );
  INV_X4 u4_sll_454_U14 ( .A(u4_sll_454_n22), .ZN(u4_sll_454_n20) );
  INV_X4 u4_sll_454_U13 ( .A(u4_sll_454_SHMAG_3_), .ZN(u4_sll_454_n24) );
  INV_X4 u4_sll_454_U12 ( .A(u4_sll_454_n24), .ZN(u4_sll_454_n22) );
  INV_X4 u4_sll_454_U11 ( .A(u4_sll_454_n34), .ZN(u4_sll_454_n29) );
  INV_X4 u4_sll_454_U10 ( .A(u4_sll_454_n48), .ZN(u4_sll_454_n46) );
  INV_X4 u4_sll_454_U9 ( .A(u4_sll_454_n49), .ZN(u4_sll_454_n45) );
  INV_X4 u4_sll_454_U8 ( .A(u4_sll_454_n34), .ZN(u4_sll_454_n30) );
  INV_X4 u4_sll_454_U7 ( .A(u4_sll_454_n33), .ZN(u4_sll_454_n31) );
  INV_X4 u4_sll_454_U6 ( .A(u4_sll_454_n33), .ZN(u4_sll_454_n32) );
  INV_X4 u4_sll_454_U5 ( .A(u4_sll_454_temp_int_SH_5_), .ZN(u4_sll_454_n51) );
  INV_X4 u4_sll_454_U4 ( .A(u4_sll_454_SHMAG_4_), .ZN(u4_sll_454_n36) );
  INV_X4 u4_sll_454_U3 ( .A(u4_sll_454_n22), .ZN(u4_sll_454_n21) );
  MUX2_X2 u4_sll_454_M1_0_1 ( .A(n6344), .B(n6446), .S(u4_sll_454_n6), .Z(
        u4_sll_454_ML_int_1__1_) );
  MUX2_X2 u4_sll_454_M1_0_2 ( .A(n6345), .B(n6344), .S(u4_sll_454_n6), .Z(
        u4_sll_454_ML_int_1__2_) );
  MUX2_X2 u4_sll_454_M1_0_3 ( .A(n6346), .B(n6345), .S(u4_sll_454_n6), .Z(
        u4_sll_454_ML_int_1__3_) );
  MUX2_X2 u4_sll_454_M1_0_4 ( .A(n6347), .B(n6346), .S(u4_sll_454_n6), .Z(
        u4_sll_454_ML_int_1__4_) );
  MUX2_X2 u4_sll_454_M1_0_5 ( .A(n6348), .B(n6347), .S(u4_sll_454_n6), .Z(
        u4_sll_454_ML_int_1__5_) );
  MUX2_X2 u4_sll_454_M1_0_6 ( .A(n6349), .B(n6348), .S(u4_sll_454_n6), .Z(
        u4_sll_454_ML_int_1__6_) );
  MUX2_X2 u4_sll_454_M1_0_7 ( .A(n6350), .B(n6349), .S(u4_sll_454_n6), .Z(
        u4_sll_454_ML_int_1__7_) );
  MUX2_X2 u4_sll_454_M1_0_8 ( .A(n6351), .B(n6350), .S(u4_sll_454_n6), .Z(
        u4_sll_454_ML_int_1__8_) );
  MUX2_X2 u4_sll_454_M1_0_9 ( .A(n6444), .B(n6351), .S(u4_sll_454_n6), .Z(
        u4_sll_454_ML_int_1__9_) );
  MUX2_X2 u4_sll_454_M1_0_10 ( .A(n6443), .B(n6444), .S(u4_sll_454_n7), .Z(
        u4_sll_454_ML_int_1__10_) );
  MUX2_X2 u4_sll_454_M1_0_11 ( .A(n6411), .B(n6443), .S(u4_sll_454_n6), .Z(
        u4_sll_454_ML_int_1__11_) );
  MUX2_X2 u4_sll_454_M1_0_12 ( .A(n6413), .B(n6411), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__12_) );
  MUX2_X2 u4_sll_454_M1_0_13 ( .A(n6414), .B(n6413), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__13_) );
  MUX2_X2 u4_sll_454_M1_0_14 ( .A(n6415), .B(n6414), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__14_) );
  MUX2_X2 u4_sll_454_M1_0_15 ( .A(n6418), .B(n6415), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__15_) );
  MUX2_X2 u4_sll_454_M1_0_16 ( .A(n6416), .B(n6418), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__16_) );
  MUX2_X2 u4_sll_454_M1_0_17 ( .A(n6417), .B(n6416), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__17_) );
  MUX2_X2 u4_sll_454_M1_0_18 ( .A(n6442), .B(n6417), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__18_) );
  MUX2_X2 u4_sll_454_M1_0_19 ( .A(n6419), .B(n6442), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__19_) );
  MUX2_X2 u4_sll_454_M1_0_20 ( .A(n6420), .B(n6419), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__20_) );
  MUX2_X2 u4_sll_454_M1_0_21 ( .A(n6421), .B(n6420), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__21_) );
  MUX2_X2 u4_sll_454_M1_0_22 ( .A(n6422), .B(n6421), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__22_) );
  MUX2_X2 u4_sll_454_M1_0_23 ( .A(n6425), .B(n6422), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__23_) );
  MUX2_X2 u4_sll_454_M1_0_24 ( .A(n6423), .B(n6425), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__24_) );
  MUX2_X2 u4_sll_454_M1_0_25 ( .A(n6424), .B(n6423), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__25_) );
  MUX2_X2 u4_sll_454_M1_0_26 ( .A(n6441), .B(n6424), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__26_) );
  MUX2_X2 u4_sll_454_M1_0_27 ( .A(n6426), .B(n6441), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__27_) );
  MUX2_X2 u4_sll_454_M1_0_28 ( .A(n6427), .B(n6426), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__28_) );
  MUX2_X2 u4_sll_454_M1_0_29 ( .A(n6428), .B(n6427), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__29_) );
  MUX2_X2 u4_sll_454_M1_0_30 ( .A(n6429), .B(n6428), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__30_) );
  MUX2_X2 u4_sll_454_M1_0_31 ( .A(n6432), .B(n6429), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__31_) );
  MUX2_X2 u4_sll_454_M1_0_32 ( .A(n6430), .B(n6432), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__32_) );
  MUX2_X2 u4_sll_454_M1_0_33 ( .A(n6431), .B(n6430), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__33_) );
  MUX2_X2 u4_sll_454_M1_0_34 ( .A(n6440), .B(n6431), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__34_) );
  MUX2_X2 u4_sll_454_M1_0_35 ( .A(n6433), .B(n6440), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__35_) );
  MUX2_X2 u4_sll_454_M1_0_36 ( .A(n6434), .B(n6433), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__36_) );
  MUX2_X2 u4_sll_454_M1_0_37 ( .A(n6435), .B(n6434), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__37_) );
  MUX2_X2 u4_sll_454_M1_0_38 ( .A(n6436), .B(n6435), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__38_) );
  MUX2_X2 u4_sll_454_M1_0_39 ( .A(n6439), .B(n6436), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__39_) );
  MUX2_X2 u4_sll_454_M1_0_40 ( .A(n6437), .B(n6439), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__40_) );
  MUX2_X2 u4_sll_454_M1_0_41 ( .A(n6438), .B(n6437), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__41_) );
  MUX2_X2 u4_sll_454_M1_0_42 ( .A(n6445), .B(n6438), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__42_) );
  MUX2_X2 u4_sll_454_M1_0_43 ( .A(n6405), .B(n6445), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__43_) );
  MUX2_X2 u4_sll_454_M1_0_44 ( .A(n6406), .B(n6405), .S(u4_sll_454_n9), .Z(
        u4_sll_454_ML_int_1__44_) );
  MUX2_X2 u4_sll_454_M1_0_45 ( .A(n6407), .B(n6406), .S(u4_sll_454_n7), .Z(
        u4_sll_454_ML_int_1__45_) );
  MUX2_X2 u4_sll_454_M1_0_46 ( .A(n6408), .B(n6407), .S(u4_sll_454_n7), .Z(
        u4_sll_454_ML_int_1__46_) );
  MUX2_X2 u4_sll_454_M1_0_47 ( .A(n6410), .B(n6408), .S(u4_sll_454_n7), .Z(
        u4_sll_454_ML_int_1__47_) );
  MUX2_X2 u4_sll_454_M1_0_48 ( .A(n6409), .B(n6410), .S(u4_sll_454_n7), .Z(
        u4_sll_454_ML_int_1__48_) );
  MUX2_X2 u4_sll_454_M1_0_49 ( .A(n6367), .B(n6409), .S(u4_sll_454_n7), .Z(
        u4_sll_454_ML_int_1__49_) );
  MUX2_X2 u4_sll_454_M1_0_50 ( .A(fract_denorm[50]), .B(n6367), .S(
        u4_sll_454_n7), .Z(u4_sll_454_ML_int_1__50_) );
  MUX2_X2 u4_sll_454_M1_0_51 ( .A(fract_denorm[51]), .B(fract_denorm[50]), .S(
        u4_sll_454_n7), .Z(u4_sll_454_ML_int_1__51_) );
  MUX2_X2 u4_sll_454_M1_0_52 ( .A(fract_denorm[52]), .B(fract_denorm[51]), .S(
        u4_sll_454_n7), .Z(u4_sll_454_ML_int_1__52_) );
  MUX2_X2 u4_sll_454_M1_0_53 ( .A(fract_denorm[53]), .B(fract_denorm[52]), .S(
        u4_sll_454_n7), .Z(u4_sll_454_ML_int_1__53_) );
  MUX2_X2 u4_sll_454_M1_0_54 ( .A(fract_denorm[54]), .B(fract_denorm[53]), .S(
        u4_sll_454_n7), .Z(u4_sll_454_ML_int_1__54_) );
  MUX2_X2 u4_sll_454_M1_0_55 ( .A(fract_denorm[55]), .B(fract_denorm[54]), .S(
        u4_sll_454_n7), .Z(u4_sll_454_ML_int_1__55_) );
  MUX2_X2 u4_sll_454_M1_0_56 ( .A(fract_denorm[56]), .B(fract_denorm[55]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__56_) );
  MUX2_X2 u4_sll_454_M1_0_57 ( .A(fract_denorm[57]), .B(fract_denorm[56]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__57_) );
  MUX2_X2 u4_sll_454_M1_0_58 ( .A(fract_denorm[58]), .B(fract_denorm[57]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__58_) );
  MUX2_X2 u4_sll_454_M1_0_59 ( .A(fract_denorm[59]), .B(fract_denorm[58]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__59_) );
  MUX2_X2 u4_sll_454_M1_0_60 ( .A(fract_denorm[60]), .B(fract_denorm[59]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__60_) );
  MUX2_X2 u4_sll_454_M1_0_61 ( .A(fract_denorm[61]), .B(fract_denorm[60]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__61_) );
  MUX2_X2 u4_sll_454_M1_0_62 ( .A(fract_denorm[62]), .B(fract_denorm[61]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__62_) );
  MUX2_X2 u4_sll_454_M1_0_63 ( .A(fract_denorm[63]), .B(fract_denorm[62]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__63_) );
  MUX2_X2 u4_sll_454_M1_0_64 ( .A(fract_denorm[64]), .B(fract_denorm[63]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__64_) );
  MUX2_X2 u4_sll_454_M1_0_65 ( .A(fract_denorm[65]), .B(fract_denorm[64]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__65_) );
  MUX2_X2 u4_sll_454_M1_0_66 ( .A(fract_denorm[66]), .B(fract_denorm[65]), .S(
        u4_sll_454_n7), .Z(u4_sll_454_ML_int_1__66_) );
  MUX2_X2 u4_sll_454_M1_0_67 ( .A(fract_denorm[67]), .B(fract_denorm[66]), .S(
        u4_sll_454_n9), .Z(u4_sll_454_ML_int_1__67_) );
  MUX2_X2 u4_sll_454_M1_0_68 ( .A(fract_denorm[68]), .B(fract_denorm[67]), .S(
        u4_sll_454_n9), .Z(u4_sll_454_ML_int_1__68_) );
  MUX2_X2 u4_sll_454_M1_0_69 ( .A(fract_denorm[69]), .B(fract_denorm[68]), .S(
        u4_sll_454_n9), .Z(u4_sll_454_ML_int_1__69_) );
  MUX2_X2 u4_sll_454_M1_0_70 ( .A(fract_denorm[70]), .B(fract_denorm[69]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__70_) );
  MUX2_X2 u4_sll_454_M1_0_71 ( .A(fract_denorm[71]), .B(fract_denorm[70]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__71_) );
  MUX2_X2 u4_sll_454_M1_0_72 ( .A(fract_denorm[72]), .B(fract_denorm[71]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__72_) );
  MUX2_X2 u4_sll_454_M1_0_73 ( .A(fract_denorm[73]), .B(fract_denorm[72]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__73_) );
  MUX2_X2 u4_sll_454_M1_0_74 ( .A(fract_denorm[74]), .B(fract_denorm[73]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__74_) );
  MUX2_X2 u4_sll_454_M1_0_75 ( .A(fract_denorm[75]), .B(fract_denorm[74]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__75_) );
  MUX2_X2 u4_sll_454_M1_0_76 ( .A(fract_denorm[76]), .B(fract_denorm[75]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__76_) );
  MUX2_X2 u4_sll_454_M1_0_77 ( .A(fract_denorm[77]), .B(fract_denorm[76]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__77_) );
  MUX2_X2 u4_sll_454_M1_0_78 ( .A(fract_denorm[78]), .B(fract_denorm[77]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__78_) );
  MUX2_X2 u4_sll_454_M1_0_79 ( .A(fract_denorm[79]), .B(fract_denorm[78]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__79_) );
  MUX2_X2 u4_sll_454_M1_0_80 ( .A(fract_denorm[80]), .B(fract_denorm[79]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__80_) );
  MUX2_X2 u4_sll_454_M1_0_81 ( .A(fract_denorm[81]), .B(fract_denorm[80]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__81_) );
  MUX2_X2 u4_sll_454_M1_0_82 ( .A(fract_denorm[82]), .B(fract_denorm[81]), .S(
        u4_sll_454_n6), .Z(u4_sll_454_ML_int_1__82_) );
  MUX2_X2 u4_sll_454_M1_0_83 ( .A(fract_denorm[83]), .B(fract_denorm[82]), .S(
        u4_sll_454_n6), .Z(u4_sll_454_ML_int_1__83_) );
  MUX2_X2 u4_sll_454_M1_0_84 ( .A(fract_denorm[84]), .B(fract_denorm[83]), .S(
        u4_sll_454_n6), .Z(u4_sll_454_ML_int_1__84_) );
  MUX2_X2 u4_sll_454_M1_0_85 ( .A(fract_denorm[85]), .B(fract_denorm[84]), .S(
        u4_sll_454_n6), .Z(u4_sll_454_ML_int_1__85_) );
  MUX2_X2 u4_sll_454_M1_0_86 ( .A(fract_denorm[86]), .B(fract_denorm[85]), .S(
        u4_sll_454_n6), .Z(u4_sll_454_ML_int_1__86_) );
  MUX2_X2 u4_sll_454_M1_0_87 ( .A(fract_denorm[87]), .B(fract_denorm[86]), .S(
        u4_sll_454_n6), .Z(u4_sll_454_ML_int_1__87_) );
  MUX2_X2 u4_sll_454_M1_0_88 ( .A(fract_denorm[88]), .B(fract_denorm[87]), .S(
        u4_sll_454_n6), .Z(u4_sll_454_ML_int_1__88_) );
  MUX2_X2 u4_sll_454_M1_0_89 ( .A(fract_denorm[89]), .B(fract_denorm[88]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__89_) );
  MUX2_X2 u4_sll_454_M1_0_90 ( .A(fract_denorm[90]), .B(fract_denorm[89]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__90_) );
  MUX2_X2 u4_sll_454_M1_0_91 ( .A(fract_denorm[91]), .B(fract_denorm[90]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__91_) );
  MUX2_X2 u4_sll_454_M1_0_92 ( .A(fract_denorm[92]), .B(fract_denorm[91]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__92_) );
  MUX2_X2 u4_sll_454_M1_0_93 ( .A(fract_denorm[93]), .B(fract_denorm[92]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__93_) );
  MUX2_X2 u4_sll_454_M1_0_94 ( .A(fract_denorm[94]), .B(fract_denorm[93]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__94_) );
  MUX2_X2 u4_sll_454_M1_0_95 ( .A(fract_denorm[95]), .B(fract_denorm[94]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__95_) );
  MUX2_X2 u4_sll_454_M1_0_96 ( .A(fract_denorm[96]), .B(fract_denorm[95]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__96_) );
  MUX2_X2 u4_sll_454_M1_0_97 ( .A(fract_denorm[97]), .B(fract_denorm[96]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__97_) );
  MUX2_X2 u4_sll_454_M1_0_98 ( .A(fract_denorm[98]), .B(fract_denorm[97]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__98_) );
  MUX2_X2 u4_sll_454_M1_0_99 ( .A(fract_denorm[99]), .B(fract_denorm[98]), .S(
        u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__99_) );
  MUX2_X2 u4_sll_454_M1_0_100 ( .A(fract_denorm[100]), .B(fract_denorm[99]), 
        .S(u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__100_) );
  MUX2_X2 u4_sll_454_M1_0_101 ( .A(fract_denorm[101]), .B(fract_denorm[100]), 
        .S(u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__101_) );
  MUX2_X2 u4_sll_454_M1_0_102 ( .A(fract_denorm[102]), .B(fract_denorm[101]), 
        .S(u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__102_) );
  MUX2_X2 u4_sll_454_M1_0_103 ( .A(fract_denorm[103]), .B(fract_denorm[102]), 
        .S(u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__103_) );
  MUX2_X2 u4_sll_454_M1_0_104 ( .A(fract_denorm[104]), .B(fract_denorm[103]), 
        .S(u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__104_) );
  MUX2_X2 u4_sll_454_M1_0_105 ( .A(fract_denorm[105]), .B(fract_denorm[104]), 
        .S(u4_sll_454_n8), .Z(u4_sll_454_ML_int_1__105_) );
  MUX2_X2 u4_sll_454_M1_1_2 ( .A(u4_sll_454_ML_int_1__2_), .B(
        u4_sll_454_ML_int_1__0_), .S(u4_sll_454_n10), .Z(
        u4_sll_454_ML_int_2__2_) );
  MUX2_X2 u4_sll_454_M1_1_3 ( .A(u4_sll_454_ML_int_1__3_), .B(
        u4_sll_454_ML_int_1__1_), .S(u4_sll_454_n10), .Z(
        u4_sll_454_ML_int_2__3_) );
  MUX2_X2 u4_sll_454_M1_1_4 ( .A(u4_sll_454_ML_int_1__4_), .B(
        u4_sll_454_ML_int_1__2_), .S(u4_sll_454_n12), .Z(
        u4_sll_454_ML_int_2__4_) );
  MUX2_X2 u4_sll_454_M1_1_5 ( .A(u4_sll_454_ML_int_1__5_), .B(
        u4_sll_454_ML_int_1__3_), .S(u4_sll_454_n12), .Z(
        u4_sll_454_ML_int_2__5_) );
  MUX2_X2 u4_sll_454_M1_1_6 ( .A(u4_sll_454_ML_int_1__6_), .B(
        u4_sll_454_ML_int_1__4_), .S(u4_sll_454_n10), .Z(
        u4_sll_454_ML_int_2__6_) );
  MUX2_X2 u4_sll_454_M1_1_7 ( .A(u4_sll_454_ML_int_1__7_), .B(
        u4_sll_454_ML_int_1__5_), .S(u4_sll_454_n10), .Z(
        u4_sll_454_ML_int_2__7_) );
  MUX2_X2 u4_sll_454_M1_1_8 ( .A(u4_sll_454_ML_int_1__8_), .B(
        u4_sll_454_ML_int_1__6_), .S(u4_sll_454_n12), .Z(
        u4_sll_454_ML_int_2__8_) );
  MUX2_X2 u4_sll_454_M1_1_9 ( .A(u4_sll_454_ML_int_1__9_), .B(
        u4_sll_454_ML_int_1__7_), .S(u4_sll_454_n12), .Z(
        u4_sll_454_ML_int_2__9_) );
  MUX2_X2 u4_sll_454_M1_1_10 ( .A(u4_sll_454_ML_int_1__10_), .B(
        u4_sll_454_ML_int_1__8_), .S(u4_sll_454_n12), .Z(
        u4_sll_454_ML_int_2__10_) );
  MUX2_X2 u4_sll_454_M1_1_11 ( .A(u4_sll_454_ML_int_1__11_), .B(
        u4_sll_454_ML_int_1__9_), .S(u4_sll_454_n10), .Z(
        u4_sll_454_ML_int_2__11_) );
  MUX2_X2 u4_sll_454_M1_1_12 ( .A(u4_sll_454_ML_int_1__12_), .B(
        u4_sll_454_ML_int_1__10_), .S(u4_sll_454_n10), .Z(
        u4_sll_454_ML_int_2__12_) );
  MUX2_X2 u4_sll_454_M1_1_13 ( .A(u4_sll_454_ML_int_1__13_), .B(
        u4_sll_454_ML_int_1__11_), .S(u4_sll_454_n12), .Z(
        u4_sll_454_ML_int_2__13_) );
  MUX2_X2 u4_sll_454_M1_1_14 ( .A(u4_sll_454_ML_int_1__14_), .B(
        u4_sll_454_ML_int_1__12_), .S(u4_sll_454_n12), .Z(
        u4_sll_454_ML_int_2__14_) );
  MUX2_X2 u4_sll_454_M1_1_15 ( .A(u4_sll_454_ML_int_1__15_), .B(
        u4_sll_454_ML_int_1__13_), .S(u4_sll_454_n12), .Z(
        u4_sll_454_ML_int_2__15_) );
  MUX2_X2 u4_sll_454_M1_1_16 ( .A(u4_sll_454_ML_int_1__16_), .B(
        u4_sll_454_ML_int_1__14_), .S(u4_sll_454_n12), .Z(
        u4_sll_454_ML_int_2__16_) );
  MUX2_X2 u4_sll_454_M1_1_17 ( .A(u4_sll_454_ML_int_1__17_), .B(
        u4_sll_454_ML_int_1__15_), .S(u4_sll_454_n12), .Z(
        u4_sll_454_ML_int_2__17_) );
  MUX2_X2 u4_sll_454_M1_1_18 ( .A(u4_sll_454_ML_int_1__18_), .B(
        u4_sll_454_ML_int_1__16_), .S(u4_sll_454_n12), .Z(
        u4_sll_454_ML_int_2__18_) );
  MUX2_X2 u4_sll_454_M1_1_19 ( .A(u4_sll_454_ML_int_1__19_), .B(
        u4_sll_454_ML_int_1__17_), .S(u4_sll_454_n12), .Z(
        u4_sll_454_ML_int_2__19_) );
  MUX2_X2 u4_sll_454_M1_1_20 ( .A(u4_sll_454_ML_int_1__20_), .B(
        u4_sll_454_ML_int_1__18_), .S(u4_sll_454_n12), .Z(
        u4_sll_454_ML_int_2__20_) );
  MUX2_X2 u4_sll_454_M1_1_21 ( .A(u4_sll_454_ML_int_1__21_), .B(
        u4_sll_454_ML_int_1__19_), .S(u4_sll_454_n12), .Z(
        u4_sll_454_ML_int_2__21_) );
  MUX2_X2 u4_sll_454_M1_1_22 ( .A(u4_sll_454_ML_int_1__22_), .B(
        u4_sll_454_ML_int_1__20_), .S(u4_sll_454_n12), .Z(
        u4_sll_454_ML_int_2__22_) );
  MUX2_X2 u4_sll_454_M1_1_23 ( .A(u4_sll_454_ML_int_1__23_), .B(
        u4_sll_454_ML_int_1__21_), .S(u4_sll_454_n12), .Z(
        u4_sll_454_ML_int_2__23_) );
  MUX2_X2 u4_sll_454_M1_1_24 ( .A(u4_sll_454_ML_int_1__24_), .B(
        u4_sll_454_ML_int_1__22_), .S(u4_sll_454_n13), .Z(
        u4_sll_454_ML_int_2__24_) );
  MUX2_X2 u4_sll_454_M1_1_25 ( .A(u4_sll_454_ML_int_1__25_), .B(
        u4_sll_454_ML_int_1__23_), .S(u4_sll_454_n13), .Z(
        u4_sll_454_ML_int_2__25_) );
  MUX2_X2 u4_sll_454_M1_1_26 ( .A(u4_sll_454_ML_int_1__26_), .B(
        u4_sll_454_ML_int_1__24_), .S(u4_sll_454_n13), .Z(
        u4_sll_454_ML_int_2__26_) );
  MUX2_X2 u4_sll_454_M1_1_27 ( .A(u4_sll_454_ML_int_1__27_), .B(
        u4_sll_454_ML_int_1__25_), .S(u4_sll_454_n13), .Z(
        u4_sll_454_ML_int_2__27_) );
  MUX2_X2 u4_sll_454_M1_1_28 ( .A(u4_sll_454_ML_int_1__28_), .B(
        u4_sll_454_ML_int_1__26_), .S(u4_sll_454_n13), .Z(
        u4_sll_454_ML_int_2__28_) );
  MUX2_X2 u4_sll_454_M1_1_29 ( .A(u4_sll_454_ML_int_1__29_), .B(
        u4_sll_454_ML_int_1__27_), .S(u4_sll_454_n13), .Z(
        u4_sll_454_ML_int_2__29_) );
  MUX2_X2 u4_sll_454_M1_1_30 ( .A(u4_sll_454_ML_int_1__30_), .B(
        u4_sll_454_ML_int_1__28_), .S(u4_sll_454_n13), .Z(
        u4_sll_454_ML_int_2__30_) );
  MUX2_X2 u4_sll_454_M1_1_31 ( .A(u4_sll_454_ML_int_1__31_), .B(
        u4_sll_454_ML_int_1__29_), .S(u4_sll_454_n12), .Z(
        u4_sll_454_ML_int_2__31_) );
  MUX2_X2 u4_sll_454_M1_1_32 ( .A(u4_sll_454_ML_int_1__32_), .B(
        u4_sll_454_ML_int_1__30_), .S(u4_sll_454_n12), .Z(
        u4_sll_454_ML_int_2__32_) );
  MUX2_X2 u4_sll_454_M1_1_33 ( .A(u4_sll_454_ML_int_1__33_), .B(
        u4_sll_454_ML_int_1__31_), .S(u4_sll_454_n12), .Z(
        u4_sll_454_ML_int_2__33_) );
  MUX2_X2 u4_sll_454_M1_1_34 ( .A(u4_sll_454_ML_int_1__34_), .B(
        u4_sll_454_ML_int_1__32_), .S(u4_sll_454_n12), .Z(
        u4_sll_454_ML_int_2__34_) );
  MUX2_X2 u4_sll_454_M1_1_35 ( .A(u4_sll_454_ML_int_1__35_), .B(
        u4_sll_454_ML_int_1__33_), .S(u4_sll_454_n13), .Z(
        u4_sll_454_ML_int_2__35_) );
  MUX2_X2 u4_sll_454_M1_1_36 ( .A(u4_sll_454_ML_int_1__36_), .B(
        u4_sll_454_ML_int_1__34_), .S(u4_sll_454_n13), .Z(
        u4_sll_454_ML_int_2__36_) );
  MUX2_X2 u4_sll_454_M1_1_37 ( .A(u4_sll_454_ML_int_1__37_), .B(
        u4_sll_454_ML_int_1__35_), .S(u4_sll_454_n13), .Z(
        u4_sll_454_ML_int_2__37_) );
  MUX2_X2 u4_sll_454_M1_1_38 ( .A(u4_sll_454_ML_int_1__38_), .B(
        u4_sll_454_ML_int_1__36_), .S(u4_sll_454_n13), .Z(
        u4_sll_454_ML_int_2__38_) );
  MUX2_X2 u4_sll_454_M1_1_39 ( .A(u4_sll_454_ML_int_1__39_), .B(
        u4_sll_454_ML_int_1__37_), .S(u4_sll_454_n13), .Z(
        u4_sll_454_ML_int_2__39_) );
  MUX2_X2 u4_sll_454_M1_1_40 ( .A(u4_sll_454_ML_int_1__40_), .B(
        u4_sll_454_ML_int_1__38_), .S(u4_sll_454_n13), .Z(
        u4_sll_454_ML_int_2__40_) );
  MUX2_X2 u4_sll_454_M1_1_41 ( .A(u4_sll_454_ML_int_1__41_), .B(
        u4_sll_454_ML_int_1__39_), .S(u4_sll_454_n13), .Z(
        u4_sll_454_ML_int_2__41_) );
  MUX2_X2 u4_sll_454_M1_1_42 ( .A(u4_sll_454_ML_int_1__42_), .B(
        u4_sll_454_ML_int_1__40_), .S(u4_sll_454_n13), .Z(
        u4_sll_454_ML_int_2__42_) );
  MUX2_X2 u4_sll_454_M1_1_43 ( .A(u4_sll_454_ML_int_1__43_), .B(
        u4_sll_454_ML_int_1__41_), .S(u4_sll_454_n13), .Z(
        u4_sll_454_ML_int_2__43_) );
  MUX2_X2 u4_sll_454_M1_1_44 ( .A(u4_sll_454_ML_int_1__44_), .B(
        u4_sll_454_ML_int_1__42_), .S(u4_sll_454_n13), .Z(
        u4_sll_454_ML_int_2__44_) );
  MUX2_X2 u4_sll_454_M1_1_45 ( .A(u4_sll_454_ML_int_1__45_), .B(
        u4_sll_454_ML_int_1__43_), .S(u4_sll_454_n13), .Z(
        u4_sll_454_ML_int_2__45_) );
  MUX2_X2 u4_sll_454_M1_1_46 ( .A(u4_sll_454_ML_int_1__46_), .B(
        u4_sll_454_ML_int_1__44_), .S(u4_sll_454_n10), .Z(
        u4_sll_454_ML_int_2__46_) );
  MUX2_X2 u4_sll_454_M1_1_47 ( .A(u4_sll_454_ML_int_1__47_), .B(
        u4_sll_454_ML_int_1__45_), .S(u4_sll_454_n10), .Z(
        u4_sll_454_ML_int_2__47_) );
  MUX2_X2 u4_sll_454_M1_1_48 ( .A(u4_sll_454_ML_int_1__48_), .B(
        u4_sll_454_ML_int_1__46_), .S(u4_sll_454_n10), .Z(
        u4_sll_454_ML_int_2__48_) );
  MUX2_X2 u4_sll_454_M1_1_49 ( .A(u4_sll_454_ML_int_1__49_), .B(
        u4_sll_454_ML_int_1__47_), .S(u4_sll_454_n10), .Z(
        u4_sll_454_ML_int_2__49_) );
  MUX2_X2 u4_sll_454_M1_1_50 ( .A(u4_sll_454_ML_int_1__50_), .B(
        u4_sll_454_ML_int_1__48_), .S(u4_sll_454_n10), .Z(
        u4_sll_454_ML_int_2__50_) );
  MUX2_X2 u4_sll_454_M1_1_51 ( .A(u4_sll_454_ML_int_1__51_), .B(
        u4_sll_454_ML_int_1__49_), .S(u4_sll_454_n10), .Z(
        u4_sll_454_ML_int_2__51_) );
  MUX2_X2 u4_sll_454_M1_1_52 ( .A(u4_sll_454_ML_int_1__52_), .B(
        u4_sll_454_ML_int_1__50_), .S(u4_sll_454_n10), .Z(
        u4_sll_454_ML_int_2__52_) );
  MUX2_X2 u4_sll_454_M1_1_53 ( .A(u4_sll_454_ML_int_1__53_), .B(
        u4_sll_454_ML_int_1__51_), .S(u4_sll_454_n10), .Z(
        u4_sll_454_ML_int_2__53_) );
  MUX2_X2 u4_sll_454_M1_1_54 ( .A(u4_sll_454_ML_int_1__54_), .B(
        u4_sll_454_ML_int_1__52_), .S(u4_sll_454_n10), .Z(
        u4_sll_454_ML_int_2__54_) );
  MUX2_X2 u4_sll_454_M1_1_55 ( .A(u4_sll_454_ML_int_1__55_), .B(
        u4_sll_454_ML_int_1__53_), .S(u4_sll_454_n10), .Z(
        u4_sll_454_ML_int_2__55_) );
  MUX2_X2 u4_sll_454_M1_1_56 ( .A(u4_sll_454_ML_int_1__56_), .B(
        u4_sll_454_ML_int_1__54_), .S(u4_sll_454_n10), .Z(
        u4_sll_454_ML_int_2__56_) );
  MUX2_X2 u4_sll_454_M1_1_57 ( .A(u4_sll_454_ML_int_1__57_), .B(
        u4_sll_454_ML_int_1__55_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__57_) );
  MUX2_X2 u4_sll_454_M1_1_58 ( .A(u4_sll_454_ML_int_1__58_), .B(
        u4_sll_454_ML_int_1__56_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__58_) );
  MUX2_X2 u4_sll_454_M1_1_59 ( .A(u4_sll_454_ML_int_1__59_), .B(
        u4_sll_454_ML_int_1__57_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__59_) );
  MUX2_X2 u4_sll_454_M1_1_60 ( .A(u4_sll_454_ML_int_1__60_), .B(
        u4_sll_454_ML_int_1__58_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__60_) );
  MUX2_X2 u4_sll_454_M1_1_61 ( .A(u4_sll_454_ML_int_1__61_), .B(
        u4_sll_454_ML_int_1__59_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__61_) );
  MUX2_X2 u4_sll_454_M1_1_62 ( .A(u4_sll_454_ML_int_1__62_), .B(
        u4_sll_454_ML_int_1__60_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__62_) );
  MUX2_X2 u4_sll_454_M1_1_63 ( .A(u4_sll_454_ML_int_1__63_), .B(
        u4_sll_454_ML_int_1__61_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__63_) );
  MUX2_X2 u4_sll_454_M1_1_64 ( .A(u4_sll_454_ML_int_1__64_), .B(
        u4_sll_454_ML_int_1__62_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__64_) );
  MUX2_X2 u4_sll_454_M1_1_65 ( .A(u4_sll_454_ML_int_1__65_), .B(
        u4_sll_454_ML_int_1__63_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__65_) );
  MUX2_X2 u4_sll_454_M1_1_66 ( .A(u4_sll_454_ML_int_1__66_), .B(
        u4_sll_454_ML_int_1__64_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__66_) );
  MUX2_X2 u4_sll_454_M1_1_67 ( .A(u4_sll_454_ML_int_1__67_), .B(
        u4_sll_454_ML_int_1__65_), .S(u4_sll_454_n10), .Z(
        u4_sll_454_ML_int_2__67_) );
  MUX2_X2 u4_sll_454_M1_1_68 ( .A(u4_sll_454_ML_int_1__68_), .B(
        u4_sll_454_ML_int_1__66_), .S(u4_sll_454_n12), .Z(
        u4_sll_454_ML_int_2__68_) );
  MUX2_X2 u4_sll_454_M1_1_69 ( .A(u4_sll_454_ML_int_1__69_), .B(
        u4_sll_454_ML_int_1__67_), .S(u4_sll_454_n12), .Z(
        u4_sll_454_ML_int_2__69_) );
  MUX2_X2 u4_sll_454_M1_1_70 ( .A(u4_sll_454_ML_int_1__70_), .B(
        u4_sll_454_ML_int_1__68_), .S(u4_sll_454_n12), .Z(
        u4_sll_454_ML_int_2__70_) );
  MUX2_X2 u4_sll_454_M1_1_71 ( .A(u4_sll_454_ML_int_1__71_), .B(
        u4_sll_454_ML_int_1__69_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__71_) );
  MUX2_X2 u4_sll_454_M1_1_72 ( .A(u4_sll_454_ML_int_1__72_), .B(
        u4_sll_454_ML_int_1__70_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__72_) );
  MUX2_X2 u4_sll_454_M1_1_73 ( .A(u4_sll_454_ML_int_1__73_), .B(
        u4_sll_454_ML_int_1__71_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__73_) );
  MUX2_X2 u4_sll_454_M1_1_74 ( .A(u4_sll_454_ML_int_1__74_), .B(
        u4_sll_454_ML_int_1__72_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__74_) );
  MUX2_X2 u4_sll_454_M1_1_75 ( .A(u4_sll_454_ML_int_1__75_), .B(
        u4_sll_454_ML_int_1__73_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__75_) );
  MUX2_X2 u4_sll_454_M1_1_76 ( .A(u4_sll_454_ML_int_1__76_), .B(
        u4_sll_454_ML_int_1__74_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__76_) );
  MUX2_X2 u4_sll_454_M1_1_77 ( .A(u4_sll_454_ML_int_1__77_), .B(
        u4_sll_454_ML_int_1__75_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__77_) );
  MUX2_X2 u4_sll_454_M1_1_78 ( .A(u4_sll_454_ML_int_1__78_), .B(
        u4_sll_454_ML_int_1__76_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__78_) );
  MUX2_X2 u4_sll_454_M1_1_79 ( .A(u4_sll_454_ML_int_1__79_), .B(
        u4_sll_454_ML_int_1__77_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__79_) );
  MUX2_X2 u4_sll_454_M1_1_80 ( .A(u4_sll_454_ML_int_1__80_), .B(
        u4_sll_454_ML_int_1__78_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__80_) );
  MUX2_X2 u4_sll_454_M1_1_81 ( .A(u4_sll_454_ML_int_1__81_), .B(
        u4_sll_454_ML_int_1__79_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__81_) );
  MUX2_X2 u4_sll_454_M1_1_82 ( .A(u4_sll_454_ML_int_1__82_), .B(
        u4_sll_454_ML_int_1__80_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__82_) );
  MUX2_X2 u4_sll_454_M1_1_83 ( .A(u4_sll_454_ML_int_1__83_), .B(
        u4_sll_454_ML_int_1__81_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__83_) );
  MUX2_X2 u4_sll_454_M1_1_84 ( .A(u4_sll_454_ML_int_1__84_), .B(
        u4_sll_454_ML_int_1__82_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__84_) );
  MUX2_X2 u4_sll_454_M1_1_85 ( .A(u4_sll_454_ML_int_1__85_), .B(
        u4_sll_454_ML_int_1__83_), .S(u4_sll_454_n12), .Z(
        u4_sll_454_ML_int_2__85_) );
  MUX2_X2 u4_sll_454_M1_1_86 ( .A(u4_sll_454_ML_int_1__86_), .B(
        u4_sll_454_ML_int_1__84_), .S(u4_sll_454_n13), .Z(
        u4_sll_454_ML_int_2__86_) );
  MUX2_X2 u4_sll_454_M1_1_87 ( .A(u4_sll_454_ML_int_1__87_), .B(
        u4_sll_454_ML_int_1__85_), .S(u4_sll_454_n12), .Z(
        u4_sll_454_ML_int_2__87_) );
  MUX2_X2 u4_sll_454_M1_1_88 ( .A(u4_sll_454_ML_int_1__88_), .B(
        u4_sll_454_ML_int_1__86_), .S(u4_sll_454_n13), .Z(
        u4_sll_454_ML_int_2__88_) );
  MUX2_X2 u4_sll_454_M1_1_89 ( .A(u4_sll_454_ML_int_1__89_), .B(
        u4_sll_454_ML_int_1__87_), .S(u4_sll_454_n12), .Z(
        u4_sll_454_ML_int_2__89_) );
  MUX2_X2 u4_sll_454_M1_1_90 ( .A(u4_sll_454_ML_int_1__90_), .B(
        u4_sll_454_ML_int_1__88_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__90_) );
  MUX2_X2 u4_sll_454_M1_1_91 ( .A(u4_sll_454_ML_int_1__91_), .B(
        u4_sll_454_ML_int_1__89_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__91_) );
  MUX2_X2 u4_sll_454_M1_1_92 ( .A(u4_sll_454_ML_int_1__92_), .B(
        u4_sll_454_ML_int_1__90_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__92_) );
  MUX2_X2 u4_sll_454_M1_1_93 ( .A(u4_sll_454_ML_int_1__93_), .B(
        u4_sll_454_ML_int_1__91_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__93_) );
  MUX2_X2 u4_sll_454_M1_1_94 ( .A(u4_sll_454_ML_int_1__94_), .B(
        u4_sll_454_ML_int_1__92_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__94_) );
  MUX2_X2 u4_sll_454_M1_1_95 ( .A(u4_sll_454_ML_int_1__95_), .B(
        u4_sll_454_ML_int_1__93_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__95_) );
  MUX2_X2 u4_sll_454_M1_1_96 ( .A(u4_sll_454_ML_int_1__96_), .B(
        u4_sll_454_ML_int_1__94_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__96_) );
  MUX2_X2 u4_sll_454_M1_1_97 ( .A(u4_sll_454_ML_int_1__97_), .B(
        u4_sll_454_ML_int_1__95_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__97_) );
  MUX2_X2 u4_sll_454_M1_1_98 ( .A(u4_sll_454_ML_int_1__98_), .B(
        u4_sll_454_ML_int_1__96_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__98_) );
  MUX2_X2 u4_sll_454_M1_1_99 ( .A(u4_sll_454_ML_int_1__99_), .B(
        u4_sll_454_ML_int_1__97_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__99_) );
  MUX2_X2 u4_sll_454_M1_1_100 ( .A(u4_sll_454_ML_int_1__100_), .B(
        u4_sll_454_ML_int_1__98_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__100_) );
  MUX2_X2 u4_sll_454_M1_1_101 ( .A(u4_sll_454_ML_int_1__101_), .B(
        u4_sll_454_ML_int_1__99_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__101_) );
  MUX2_X2 u4_sll_454_M1_1_102 ( .A(u4_sll_454_ML_int_1__102_), .B(
        u4_sll_454_ML_int_1__100_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__102_) );
  MUX2_X2 u4_sll_454_M1_1_103 ( .A(u4_sll_454_ML_int_1__103_), .B(
        u4_sll_454_ML_int_1__101_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__103_) );
  MUX2_X2 u4_sll_454_M1_1_104 ( .A(u4_sll_454_ML_int_1__104_), .B(
        u4_sll_454_ML_int_1__102_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__104_) );
  MUX2_X2 u4_sll_454_M1_1_105 ( .A(u4_sll_454_ML_int_1__105_), .B(
        u4_sll_454_ML_int_1__103_), .S(u4_sll_454_n11), .Z(
        u4_sll_454_ML_int_2__105_) );
  MUX2_X2 u4_sll_454_M1_2_4 ( .A(u4_sll_454_ML_int_2__4_), .B(
        u4_sll_454_ML_int_2__0_), .S(u4_sll_454_n17), .Z(
        u4_sll_454_ML_int_3__4_) );
  MUX2_X2 u4_sll_454_M1_2_5 ( .A(u4_sll_454_ML_int_2__5_), .B(
        u4_sll_454_ML_int_2__1_), .S(u4_sll_454_n17), .Z(
        u4_sll_454_ML_int_3__5_) );
  MUX2_X2 u4_sll_454_M1_2_6 ( .A(u4_sll_454_ML_int_2__6_), .B(
        u4_sll_454_ML_int_2__2_), .S(u4_sll_454_n17), .Z(
        u4_sll_454_ML_int_3__6_) );
  MUX2_X2 u4_sll_454_M1_2_7 ( .A(u4_sll_454_ML_int_2__7_), .B(
        u4_sll_454_ML_int_2__3_), .S(u4_sll_454_n17), .Z(
        u4_sll_454_ML_int_3__7_) );
  MUX2_X2 u4_sll_454_M1_2_8 ( .A(u4_sll_454_ML_int_2__8_), .B(
        u4_sll_454_ML_int_2__4_), .S(u4_sll_454_n17), .Z(
        u4_sll_454_ML_int_3__8_) );
  MUX2_X2 u4_sll_454_M1_2_9 ( .A(u4_sll_454_ML_int_2__9_), .B(
        u4_sll_454_ML_int_2__5_), .S(u4_sll_454_n17), .Z(
        u4_sll_454_ML_int_3__9_) );
  MUX2_X2 u4_sll_454_M1_2_10 ( .A(u4_sll_454_ML_int_2__10_), .B(
        u4_sll_454_ML_int_2__6_), .S(u4_sll_454_n17), .Z(
        u4_sll_454_ML_int_3__10_) );
  MUX2_X2 u4_sll_454_M1_2_11 ( .A(u4_sll_454_ML_int_2__11_), .B(
        u4_sll_454_ML_int_2__7_), .S(u4_sll_454_n17), .Z(
        u4_sll_454_ML_int_3__11_) );
  MUX2_X2 u4_sll_454_M1_2_12 ( .A(u4_sll_454_ML_int_2__12_), .B(
        u4_sll_454_ML_int_2__8_), .S(u4_sll_454_n17), .Z(
        u4_sll_454_ML_int_3__12_) );
  MUX2_X2 u4_sll_454_M1_2_13 ( .A(u4_sll_454_ML_int_2__13_), .B(
        u4_sll_454_ML_int_2__9_), .S(u4_sll_454_n17), .Z(
        u4_sll_454_ML_int_3__13_) );
  MUX2_X2 u4_sll_454_M1_2_14 ( .A(u4_sll_454_ML_int_2__14_), .B(
        u4_sll_454_ML_int_2__10_), .S(u4_sll_454_n17), .Z(
        u4_sll_454_ML_int_3__14_) );
  MUX2_X2 u4_sll_454_M1_2_15 ( .A(u4_sll_454_ML_int_2__15_), .B(
        u4_sll_454_ML_int_2__11_), .S(u4_sll_454_n14), .Z(
        u4_sll_454_ML_int_3__15_) );
  MUX2_X2 u4_sll_454_M1_2_16 ( .A(u4_sll_454_ML_int_2__16_), .B(
        u4_sll_454_ML_int_2__12_), .S(u4_sll_454_n17), .Z(
        u4_sll_454_ML_int_3__16_) );
  MUX2_X2 u4_sll_454_M1_2_17 ( .A(u4_sll_454_ML_int_2__17_), .B(
        u4_sll_454_ML_int_2__13_), .S(u4_sll_454_n17), .Z(
        u4_sll_454_ML_int_3__17_) );
  MUX2_X2 u4_sll_454_M1_2_18 ( .A(u4_sll_454_ML_int_2__18_), .B(
        u4_sll_454_ML_int_2__14_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__18_) );
  MUX2_X2 u4_sll_454_M1_2_19 ( .A(u4_sll_454_ML_int_2__19_), .B(
        u4_sll_454_ML_int_2__15_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__19_) );
  MUX2_X2 u4_sll_454_M1_2_20 ( .A(u4_sll_454_ML_int_2__20_), .B(
        u4_sll_454_ML_int_2__16_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__20_) );
  MUX2_X2 u4_sll_454_M1_2_21 ( .A(u4_sll_454_ML_int_2__21_), .B(
        u4_sll_454_ML_int_2__17_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__21_) );
  MUX2_X2 u4_sll_454_M1_2_22 ( .A(u4_sll_454_ML_int_2__22_), .B(
        u4_sll_454_ML_int_2__18_), .S(u4_sll_454_n17), .Z(
        u4_sll_454_ML_int_3__22_) );
  MUX2_X2 u4_sll_454_M1_2_23 ( .A(u4_sll_454_ML_int_2__23_), .B(
        u4_sll_454_ML_int_2__19_), .S(u4_sll_454_n14), .Z(
        u4_sll_454_ML_int_3__23_) );
  MUX2_X2 u4_sll_454_M1_2_24 ( .A(u4_sll_454_ML_int_2__24_), .B(
        u4_sll_454_ML_int_2__20_), .S(u4_sll_454_n17), .Z(
        u4_sll_454_ML_int_3__24_) );
  MUX2_X2 u4_sll_454_M1_2_25 ( .A(u4_sll_454_ML_int_2__25_), .B(
        u4_sll_454_ML_int_2__21_), .S(u4_sll_454_n16), .Z(
        u4_sll_454_ML_int_3__25_) );
  MUX2_X2 u4_sll_454_M1_2_26 ( .A(u4_sll_454_ML_int_2__26_), .B(
        u4_sll_454_ML_int_2__22_), .S(u4_sll_454_n16), .Z(
        u4_sll_454_ML_int_3__26_) );
  MUX2_X2 u4_sll_454_M1_2_27 ( .A(u4_sll_454_ML_int_2__27_), .B(
        u4_sll_454_ML_int_2__23_), .S(u4_sll_454_n16), .Z(
        u4_sll_454_ML_int_3__27_) );
  MUX2_X2 u4_sll_454_M1_2_28 ( .A(u4_sll_454_ML_int_2__28_), .B(
        u4_sll_454_ML_int_2__24_), .S(u4_sll_454_n16), .Z(
        u4_sll_454_ML_int_3__28_) );
  MUX2_X2 u4_sll_454_M1_2_29 ( .A(u4_sll_454_ML_int_2__29_), .B(
        u4_sll_454_ML_int_2__25_), .S(u4_sll_454_n16), .Z(
        u4_sll_454_ML_int_3__29_) );
  MUX2_X2 u4_sll_454_M1_2_30 ( .A(u4_sll_454_ML_int_2__30_), .B(
        u4_sll_454_ML_int_2__26_), .S(u4_sll_454_n16), .Z(
        u4_sll_454_ML_int_3__30_) );
  MUX2_X2 u4_sll_454_M1_2_31 ( .A(u4_sll_454_ML_int_2__31_), .B(
        u4_sll_454_ML_int_2__27_), .S(u4_sll_454_n16), .Z(
        u4_sll_454_ML_int_3__31_) );
  MUX2_X2 u4_sll_454_M1_2_32 ( .A(u4_sll_454_ML_int_2__32_), .B(
        u4_sll_454_ML_int_2__28_), .S(u4_sll_454_n16), .Z(
        u4_sll_454_ML_int_3__32_) );
  MUX2_X2 u4_sll_454_M1_2_33 ( .A(u4_sll_454_ML_int_2__33_), .B(
        u4_sll_454_ML_int_2__29_), .S(u4_sll_454_n17), .Z(
        u4_sll_454_ML_int_3__33_) );
  MUX2_X2 u4_sll_454_M1_2_34 ( .A(u4_sll_454_ML_int_2__34_), .B(
        u4_sll_454_ML_int_2__30_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__34_) );
  MUX2_X2 u4_sll_454_M1_2_35 ( .A(u4_sll_454_ML_int_2__35_), .B(
        u4_sll_454_ML_int_2__31_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__35_) );
  MUX2_X2 u4_sll_454_M1_2_36 ( .A(u4_sll_454_ML_int_2__36_), .B(
        u4_sll_454_ML_int_2__32_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__36_) );
  MUX2_X2 u4_sll_454_M1_2_37 ( .A(u4_sll_454_ML_int_2__37_), .B(
        u4_sll_454_ML_int_2__33_), .S(u4_sll_454_n16), .Z(
        u4_sll_454_ML_int_3__37_) );
  MUX2_X2 u4_sll_454_M1_2_38 ( .A(u4_sll_454_ML_int_2__38_), .B(
        u4_sll_454_ML_int_2__34_), .S(u4_sll_454_n16), .Z(
        u4_sll_454_ML_int_3__38_) );
  MUX2_X2 u4_sll_454_M1_2_39 ( .A(u4_sll_454_ML_int_2__39_), .B(
        u4_sll_454_ML_int_2__35_), .S(u4_sll_454_n16), .Z(
        u4_sll_454_ML_int_3__39_) );
  MUX2_X2 u4_sll_454_M1_2_40 ( .A(u4_sll_454_ML_int_2__40_), .B(
        u4_sll_454_ML_int_2__36_), .S(u4_sll_454_n16), .Z(
        u4_sll_454_ML_int_3__40_) );
  MUX2_X2 u4_sll_454_M1_2_41 ( .A(u4_sll_454_ML_int_2__41_), .B(
        u4_sll_454_ML_int_2__37_), .S(u4_sll_454_n16), .Z(
        u4_sll_454_ML_int_3__41_) );
  MUX2_X2 u4_sll_454_M1_2_42 ( .A(u4_sll_454_ML_int_2__42_), .B(
        u4_sll_454_ML_int_2__38_), .S(u4_sll_454_n16), .Z(
        u4_sll_454_ML_int_3__42_) );
  MUX2_X2 u4_sll_454_M1_2_43 ( .A(u4_sll_454_ML_int_2__43_), .B(
        u4_sll_454_ML_int_2__39_), .S(u4_sll_454_n16), .Z(
        u4_sll_454_ML_int_3__43_) );
  MUX2_X2 u4_sll_454_M1_2_44 ( .A(u4_sll_454_ML_int_2__44_), .B(
        u4_sll_454_ML_int_2__40_), .S(u4_sll_454_n16), .Z(
        u4_sll_454_ML_int_3__44_) );
  MUX2_X2 u4_sll_454_M1_2_45 ( .A(u4_sll_454_ML_int_2__45_), .B(
        u4_sll_454_ML_int_2__41_), .S(u4_sll_454_n16), .Z(
        u4_sll_454_ML_int_3__45_) );
  MUX2_X2 u4_sll_454_M1_2_46 ( .A(u4_sll_454_ML_int_2__46_), .B(
        u4_sll_454_ML_int_2__42_), .S(u4_sll_454_n16), .Z(
        u4_sll_454_ML_int_3__46_) );
  MUX2_X2 u4_sll_454_M1_2_47 ( .A(u4_sll_454_ML_int_2__47_), .B(
        u4_sll_454_ML_int_2__43_), .S(u4_sll_454_n16), .Z(
        u4_sll_454_ML_int_3__47_) );
  MUX2_X2 u4_sll_454_M1_2_48 ( .A(u4_sll_454_ML_int_2__48_), .B(
        u4_sll_454_ML_int_2__44_), .S(u4_sll_454_n14), .Z(
        u4_sll_454_ML_int_3__48_) );
  MUX2_X2 u4_sll_454_M1_2_49 ( .A(u4_sll_454_ML_int_2__49_), .B(
        u4_sll_454_ML_int_2__45_), .S(u4_sll_454_n14), .Z(
        u4_sll_454_ML_int_3__49_) );
  MUX2_X2 u4_sll_454_M1_2_50 ( .A(u4_sll_454_ML_int_2__50_), .B(
        u4_sll_454_ML_int_2__46_), .S(u4_sll_454_n14), .Z(
        u4_sll_454_ML_int_3__50_) );
  MUX2_X2 u4_sll_454_M1_2_51 ( .A(u4_sll_454_ML_int_2__51_), .B(
        u4_sll_454_ML_int_2__47_), .S(u4_sll_454_n14), .Z(
        u4_sll_454_ML_int_3__51_) );
  MUX2_X2 u4_sll_454_M1_2_52 ( .A(u4_sll_454_ML_int_2__52_), .B(
        u4_sll_454_ML_int_2__48_), .S(u4_sll_454_n14), .Z(
        u4_sll_454_ML_int_3__52_) );
  MUX2_X2 u4_sll_454_M1_2_53 ( .A(u4_sll_454_ML_int_2__53_), .B(
        u4_sll_454_ML_int_2__49_), .S(u4_sll_454_n14), .Z(
        u4_sll_454_ML_int_3__53_) );
  MUX2_X2 u4_sll_454_M1_2_54 ( .A(u4_sll_454_ML_int_2__54_), .B(
        u4_sll_454_ML_int_2__50_), .S(u4_sll_454_n14), .Z(
        u4_sll_454_ML_int_3__54_) );
  MUX2_X2 u4_sll_454_M1_2_55 ( .A(u4_sll_454_ML_int_2__55_), .B(
        u4_sll_454_ML_int_2__51_), .S(u4_sll_454_n14), .Z(
        u4_sll_454_ML_int_3__55_) );
  MUX2_X2 u4_sll_454_M1_2_56 ( .A(u4_sll_454_ML_int_2__56_), .B(
        u4_sll_454_ML_int_2__52_), .S(u4_sll_454_n14), .Z(
        u4_sll_454_ML_int_3__56_) );
  MUX2_X2 u4_sll_454_M1_2_57 ( .A(u4_sll_454_ML_int_2__57_), .B(
        u4_sll_454_ML_int_2__53_), .S(u4_sll_454_n14), .Z(
        u4_sll_454_ML_int_3__57_) );
  MUX2_X2 u4_sll_454_M1_2_58 ( .A(u4_sll_454_ML_int_2__58_), .B(
        u4_sll_454_ML_int_2__54_), .S(u4_sll_454_n14), .Z(
        u4_sll_454_ML_int_3__58_) );
  MUX2_X2 u4_sll_454_M1_2_59 ( .A(u4_sll_454_ML_int_2__59_), .B(
        u4_sll_454_ML_int_2__55_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__59_) );
  MUX2_X2 u4_sll_454_M1_2_60 ( .A(u4_sll_454_ML_int_2__60_), .B(
        u4_sll_454_ML_int_2__56_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__60_) );
  MUX2_X2 u4_sll_454_M1_2_61 ( .A(u4_sll_454_ML_int_2__61_), .B(
        u4_sll_454_ML_int_2__57_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__61_) );
  MUX2_X2 u4_sll_454_M1_2_62 ( .A(u4_sll_454_ML_int_2__62_), .B(
        u4_sll_454_ML_int_2__58_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__62_) );
  MUX2_X2 u4_sll_454_M1_2_63 ( .A(u4_sll_454_ML_int_2__63_), .B(
        u4_sll_454_ML_int_2__59_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__63_) );
  MUX2_X2 u4_sll_454_M1_2_64 ( .A(u4_sll_454_ML_int_2__64_), .B(
        u4_sll_454_ML_int_2__60_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__64_) );
  MUX2_X2 u4_sll_454_M1_2_65 ( .A(u4_sll_454_ML_int_2__65_), .B(
        u4_sll_454_ML_int_2__61_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__65_) );
  MUX2_X2 u4_sll_454_M1_2_66 ( .A(u4_sll_454_ML_int_2__66_), .B(
        u4_sll_454_ML_int_2__62_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__66_) );
  MUX2_X2 u4_sll_454_M1_2_67 ( .A(u4_sll_454_ML_int_2__67_), .B(
        u4_sll_454_ML_int_2__63_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__67_) );
  MUX2_X2 u4_sll_454_M1_2_68 ( .A(u4_sll_454_ML_int_2__68_), .B(
        u4_sll_454_ML_int_2__64_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__68_) );
  MUX2_X2 u4_sll_454_M1_2_69 ( .A(u4_sll_454_ML_int_2__69_), .B(
        u4_sll_454_ML_int_2__65_), .S(u4_sll_454_n14), .Z(
        u4_sll_454_ML_int_3__69_) );
  MUX2_X2 u4_sll_454_M1_2_70 ( .A(u4_sll_454_ML_int_2__70_), .B(
        u4_sll_454_ML_int_2__66_), .S(u4_sll_454_n14), .Z(
        u4_sll_454_ML_int_3__70_) );
  MUX2_X2 u4_sll_454_M1_2_71 ( .A(u4_sll_454_ML_int_2__71_), .B(
        u4_sll_454_ML_int_2__67_), .S(u4_sll_454_n17), .Z(
        u4_sll_454_ML_int_3__71_) );
  MUX2_X2 u4_sll_454_M1_2_72 ( .A(u4_sll_454_ML_int_2__72_), .B(
        u4_sll_454_ML_int_2__68_), .S(u4_sll_454_n16), .Z(
        u4_sll_454_ML_int_3__72_) );
  MUX2_X2 u4_sll_454_M1_2_73 ( .A(u4_sll_454_ML_int_2__73_), .B(
        u4_sll_454_ML_int_2__69_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__73_) );
  MUX2_X2 u4_sll_454_M1_2_74 ( .A(u4_sll_454_ML_int_2__74_), .B(
        u4_sll_454_ML_int_2__70_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__74_) );
  MUX2_X2 u4_sll_454_M1_2_75 ( .A(u4_sll_454_ML_int_2__75_), .B(
        u4_sll_454_ML_int_2__71_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__75_) );
  MUX2_X2 u4_sll_454_M1_2_76 ( .A(u4_sll_454_ML_int_2__76_), .B(
        u4_sll_454_ML_int_2__72_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__76_) );
  MUX2_X2 u4_sll_454_M1_2_77 ( .A(u4_sll_454_ML_int_2__77_), .B(
        u4_sll_454_ML_int_2__73_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__77_) );
  MUX2_X2 u4_sll_454_M1_2_78 ( .A(u4_sll_454_ML_int_2__78_), .B(
        u4_sll_454_ML_int_2__74_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__78_) );
  MUX2_X2 u4_sll_454_M1_2_79 ( .A(u4_sll_454_ML_int_2__79_), .B(
        u4_sll_454_ML_int_2__75_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__79_) );
  MUX2_X2 u4_sll_454_M1_2_80 ( .A(u4_sll_454_ML_int_2__80_), .B(
        u4_sll_454_ML_int_2__76_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__80_) );
  MUX2_X2 u4_sll_454_M1_2_81 ( .A(u4_sll_454_ML_int_2__81_), .B(
        u4_sll_454_ML_int_2__77_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__81_) );
  MUX2_X2 u4_sll_454_M1_2_82 ( .A(u4_sll_454_ML_int_2__82_), .B(
        u4_sll_454_ML_int_2__78_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__82_) );
  MUX2_X2 u4_sll_454_M1_2_83 ( .A(u4_sll_454_ML_int_2__83_), .B(
        u4_sll_454_ML_int_2__79_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__83_) );
  MUX2_X2 u4_sll_454_M1_2_84 ( .A(u4_sll_454_ML_int_2__84_), .B(
        u4_sll_454_ML_int_2__80_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__84_) );
  MUX2_X2 u4_sll_454_M1_2_85 ( .A(u4_sll_454_ML_int_2__85_), .B(
        u4_sll_454_ML_int_2__81_), .S(u4_sll_454_n17), .Z(
        u4_sll_454_ML_int_3__85_) );
  MUX2_X2 u4_sll_454_M1_2_86 ( .A(u4_sll_454_ML_int_2__86_), .B(
        u4_sll_454_ML_int_2__82_), .S(u4_sll_454_n17), .Z(
        u4_sll_454_ML_int_3__86_) );
  MUX2_X2 u4_sll_454_M1_2_87 ( .A(u4_sll_454_ML_int_2__87_), .B(
        u4_sll_454_ML_int_2__83_), .S(u4_sll_454_n17), .Z(
        u4_sll_454_ML_int_3__87_) );
  MUX2_X2 u4_sll_454_M1_2_88 ( .A(u4_sll_454_ML_int_2__88_), .B(
        u4_sll_454_ML_int_2__84_), .S(u4_sll_454_n17), .Z(
        u4_sll_454_ML_int_3__88_) );
  MUX2_X2 u4_sll_454_M1_2_89 ( .A(u4_sll_454_ML_int_2__89_), .B(
        u4_sll_454_ML_int_2__85_), .S(u4_sll_454_n17), .Z(
        u4_sll_454_ML_int_3__89_) );
  MUX2_X2 u4_sll_454_M1_2_90 ( .A(u4_sll_454_ML_int_2__90_), .B(
        u4_sll_454_ML_int_2__86_), .S(u4_sll_454_n17), .Z(
        u4_sll_454_ML_int_3__90_) );
  MUX2_X2 u4_sll_454_M1_2_91 ( .A(u4_sll_454_ML_int_2__91_), .B(
        u4_sll_454_ML_int_2__87_), .S(u4_sll_454_n17), .Z(
        u4_sll_454_ML_int_3__91_) );
  MUX2_X2 u4_sll_454_M1_2_92 ( .A(u4_sll_454_ML_int_2__92_), .B(
        u4_sll_454_ML_int_2__88_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__92_) );
  MUX2_X2 u4_sll_454_M1_2_93 ( .A(u4_sll_454_ML_int_2__93_), .B(
        u4_sll_454_ML_int_2__89_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__93_) );
  MUX2_X2 u4_sll_454_M1_2_94 ( .A(u4_sll_454_ML_int_2__94_), .B(
        u4_sll_454_ML_int_2__90_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__94_) );
  MUX2_X2 u4_sll_454_M1_2_95 ( .A(u4_sll_454_ML_int_2__95_), .B(
        u4_sll_454_ML_int_2__91_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__95_) );
  MUX2_X2 u4_sll_454_M1_2_96 ( .A(u4_sll_454_ML_int_2__96_), .B(
        u4_sll_454_ML_int_2__92_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__96_) );
  MUX2_X2 u4_sll_454_M1_2_97 ( .A(u4_sll_454_ML_int_2__97_), .B(
        u4_sll_454_ML_int_2__93_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__97_) );
  MUX2_X2 u4_sll_454_M1_2_98 ( .A(u4_sll_454_ML_int_2__98_), .B(
        u4_sll_454_ML_int_2__94_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__98_) );
  MUX2_X2 u4_sll_454_M1_2_99 ( .A(u4_sll_454_ML_int_2__99_), .B(
        u4_sll_454_ML_int_2__95_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__99_) );
  MUX2_X2 u4_sll_454_M1_2_100 ( .A(u4_sll_454_ML_int_2__100_), .B(
        u4_sll_454_ML_int_2__96_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__100_) );
  MUX2_X2 u4_sll_454_M1_2_101 ( .A(u4_sll_454_ML_int_2__101_), .B(
        u4_sll_454_ML_int_2__97_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__101_) );
  MUX2_X2 u4_sll_454_M1_2_102 ( .A(u4_sll_454_ML_int_2__102_), .B(
        u4_sll_454_ML_int_2__98_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__102_) );
  MUX2_X2 u4_sll_454_M1_2_103 ( .A(u4_sll_454_ML_int_2__103_), .B(
        u4_sll_454_ML_int_2__99_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__103_) );
  MUX2_X2 u4_sll_454_M1_2_104 ( .A(u4_sll_454_ML_int_2__104_), .B(
        u4_sll_454_ML_int_2__100_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__104_) );
  MUX2_X2 u4_sll_454_M1_2_105 ( .A(u4_sll_454_ML_int_2__105_), .B(
        u4_sll_454_ML_int_2__101_), .S(u4_sll_454_n15), .Z(
        u4_sll_454_ML_int_3__105_) );
  MUX2_X2 u4_sll_454_M1_3_8 ( .A(u4_sll_454_ML_int_3__8_), .B(
        u4_sll_454_ML_int_3__0_), .S(u4_sll_454_n21), .Z(
        u4_sll_454_ML_int_4__8_) );
  MUX2_X2 u4_sll_454_M1_3_9 ( .A(u4_sll_454_ML_int_3__9_), .B(
        u4_sll_454_ML_int_3__1_), .S(u4_sll_454_n21), .Z(
        u4_sll_454_ML_int_4__9_) );
  MUX2_X2 u4_sll_454_M1_3_10 ( .A(u4_sll_454_ML_int_3__10_), .B(
        u4_sll_454_ML_int_3__2_), .S(u4_sll_454_n21), .Z(
        u4_sll_454_ML_int_4__10_) );
  MUX2_X2 u4_sll_454_M1_3_11 ( .A(u4_sll_454_ML_int_3__11_), .B(
        u4_sll_454_ML_int_3__3_), .S(u4_sll_454_n21), .Z(
        u4_sll_454_ML_int_4__11_) );
  MUX2_X2 u4_sll_454_M1_3_12 ( .A(u4_sll_454_ML_int_3__12_), .B(
        u4_sll_454_ML_int_3__4_), .S(u4_sll_454_n21), .Z(
        u4_sll_454_ML_int_4__12_) );
  MUX2_X2 u4_sll_454_M1_3_13 ( .A(u4_sll_454_ML_int_3__13_), .B(
        u4_sll_454_ML_int_3__5_), .S(u4_sll_454_n21), .Z(
        u4_sll_454_ML_int_4__13_) );
  MUX2_X2 u4_sll_454_M1_3_14 ( .A(u4_sll_454_ML_int_3__14_), .B(
        u4_sll_454_ML_int_3__6_), .S(u4_sll_454_n21), .Z(
        u4_sll_454_ML_int_4__14_) );
  MUX2_X2 u4_sll_454_M1_3_15 ( .A(u4_sll_454_ML_int_3__15_), .B(
        u4_sll_454_ML_int_3__7_), .S(u4_sll_454_n21), .Z(
        u4_sll_454_ML_int_4__15_) );
  MUX2_X2 u4_sll_454_M1_3_16 ( .A(u4_sll_454_ML_int_3__16_), .B(
        u4_sll_454_ML_int_3__8_), .S(u4_sll_454_n21), .Z(
        u4_sll_454_ML_int_4__16_) );
  MUX2_X2 u4_sll_454_M1_3_17 ( .A(u4_sll_454_ML_int_3__17_), .B(
        u4_sll_454_ML_int_3__9_), .S(u4_sll_454_n21), .Z(
        u4_sll_454_ML_int_4__17_) );
  MUX2_X2 u4_sll_454_M1_3_18 ( .A(u4_sll_454_ML_int_3__18_), .B(
        u4_sll_454_ML_int_3__10_), .S(u4_sll_454_n20), .Z(
        u4_sll_454_ML_int_4__18_) );
  MUX2_X2 u4_sll_454_M1_3_19 ( .A(u4_sll_454_ML_int_3__19_), .B(
        u4_sll_454_ML_int_3__11_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__19_) );
  MUX2_X2 u4_sll_454_M1_3_20 ( .A(u4_sll_454_ML_int_3__20_), .B(
        u4_sll_454_ML_int_3__12_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__20_) );
  MUX2_X2 u4_sll_454_M1_3_21 ( .A(u4_sll_454_ML_int_3__21_), .B(
        u4_sll_454_ML_int_3__13_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__21_) );
  MUX2_X2 u4_sll_454_M1_3_22 ( .A(u4_sll_454_ML_int_3__22_), .B(
        u4_sll_454_ML_int_3__14_), .S(u4_sll_454_n21), .Z(
        u4_sll_454_ML_int_4__22_) );
  MUX2_X2 u4_sll_454_M1_3_23 ( .A(u4_sll_454_ML_int_3__23_), .B(
        u4_sll_454_ML_int_3__15_), .S(u4_sll_454_n21), .Z(
        u4_sll_454_ML_int_4__23_) );
  MUX2_X2 u4_sll_454_M1_3_24 ( .A(u4_sll_454_ML_int_3__24_), .B(
        u4_sll_454_ML_int_3__16_), .S(u4_sll_454_n21), .Z(
        u4_sll_454_ML_int_4__24_) );
  MUX2_X2 u4_sll_454_M1_3_25 ( .A(u4_sll_454_ML_int_3__25_), .B(
        u4_sll_454_ML_int_3__17_), .S(u4_sll_454_n21), .Z(
        u4_sll_454_ML_int_4__25_) );
  MUX2_X2 u4_sll_454_M1_3_26 ( .A(u4_sll_454_ML_int_3__26_), .B(
        u4_sll_454_ML_int_3__18_), .S(u4_sll_454_n21), .Z(
        u4_sll_454_ML_int_4__26_) );
  MUX2_X2 u4_sll_454_M1_3_27 ( .A(u4_sll_454_ML_int_3__27_), .B(
        u4_sll_454_ML_int_3__19_), .S(u4_sll_454_n21), .Z(
        u4_sll_454_ML_int_4__27_) );
  MUX2_X2 u4_sll_454_M1_3_28 ( .A(u4_sll_454_ML_int_3__28_), .B(
        u4_sll_454_ML_int_3__20_), .S(u4_sll_454_n21), .Z(
        u4_sll_454_ML_int_4__28_) );
  MUX2_X2 u4_sll_454_M1_3_29 ( .A(u4_sll_454_ML_int_3__29_), .B(
        u4_sll_454_ML_int_3__21_), .S(u4_sll_454_n21), .Z(
        u4_sll_454_ML_int_4__29_) );
  MUX2_X2 u4_sll_454_M1_3_30 ( .A(u4_sll_454_ML_int_3__30_), .B(
        u4_sll_454_ML_int_3__22_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__30_) );
  MUX2_X2 u4_sll_454_M1_3_31 ( .A(u4_sll_454_ML_int_3__31_), .B(
        u4_sll_454_ML_int_3__23_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__31_) );
  MUX2_X2 u4_sll_454_M1_3_32 ( .A(u4_sll_454_ML_int_3__32_), .B(
        u4_sll_454_ML_int_3__24_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__32_) );
  MUX2_X2 u4_sll_454_M1_3_33 ( .A(u4_sll_454_ML_int_3__33_), .B(
        u4_sll_454_ML_int_3__25_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__33_) );
  MUX2_X2 u4_sll_454_M1_3_34 ( .A(u4_sll_454_ML_int_3__34_), .B(
        u4_sll_454_ML_int_3__26_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__34_) );
  MUX2_X2 u4_sll_454_M1_3_35 ( .A(u4_sll_454_ML_int_3__35_), .B(
        u4_sll_454_ML_int_3__27_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__35_) );
  MUX2_X2 u4_sll_454_M1_3_36 ( .A(u4_sll_454_ML_int_3__36_), .B(
        u4_sll_454_ML_int_3__28_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__36_) );
  MUX2_X2 u4_sll_454_M1_3_37 ( .A(u4_sll_454_ML_int_3__37_), .B(
        u4_sll_454_ML_int_3__29_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__37_) );
  MUX2_X2 u4_sll_454_M1_3_38 ( .A(u4_sll_454_ML_int_3__38_), .B(
        u4_sll_454_ML_int_3__30_), .S(u4_sll_454_n24), .Z(
        u4_sll_454_ML_int_4__38_) );
  MUX2_X2 u4_sll_454_M1_3_39 ( .A(u4_sll_454_ML_int_3__39_), .B(
        u4_sll_454_ML_int_3__31_), .S(u4_sll_454_n20), .Z(
        u4_sll_454_ML_int_4__39_) );
  MUX2_X2 u4_sll_454_M1_3_40 ( .A(u4_sll_454_ML_int_3__40_), .B(
        u4_sll_454_ML_int_3__32_), .S(u4_sll_454_n19), .Z(
        u4_sll_454_ML_int_4__40_) );
  MUX2_X2 u4_sll_454_M1_3_41 ( .A(u4_sll_454_ML_int_3__41_), .B(
        u4_sll_454_ML_int_3__33_), .S(u4_sll_454_n19), .Z(
        u4_sll_454_ML_int_4__41_) );
  MUX2_X2 u4_sll_454_M1_3_42 ( .A(u4_sll_454_ML_int_3__42_), .B(
        u4_sll_454_ML_int_3__34_), .S(u4_sll_454_n19), .Z(
        u4_sll_454_ML_int_4__42_) );
  MUX2_X2 u4_sll_454_M1_3_43 ( .A(u4_sll_454_ML_int_3__43_), .B(
        u4_sll_454_ML_int_3__35_), .S(u4_sll_454_n19), .Z(
        u4_sll_454_ML_int_4__43_) );
  MUX2_X2 u4_sll_454_M1_3_44 ( .A(u4_sll_454_ML_int_3__44_), .B(
        u4_sll_454_ML_int_3__36_), .S(u4_sll_454_n19), .Z(
        u4_sll_454_ML_int_4__44_) );
  MUX2_X2 u4_sll_454_M1_3_45 ( .A(u4_sll_454_ML_int_3__45_), .B(
        u4_sll_454_ML_int_3__37_), .S(u4_sll_454_n19), .Z(
        u4_sll_454_ML_int_4__45_) );
  MUX2_X2 u4_sll_454_M1_3_46 ( .A(u4_sll_454_ML_int_3__46_), .B(
        u4_sll_454_ML_int_3__38_), .S(u4_sll_454_n19), .Z(
        u4_sll_454_ML_int_4__46_) );
  MUX2_X2 u4_sll_454_M1_3_47 ( .A(u4_sll_454_ML_int_3__47_), .B(
        u4_sll_454_ML_int_3__39_), .S(u4_sll_454_n19), .Z(
        u4_sll_454_ML_int_4__47_) );
  MUX2_X2 u4_sll_454_M1_3_48 ( .A(u4_sll_454_ML_int_3__48_), .B(
        u4_sll_454_ML_int_3__40_), .S(u4_sll_454_n19), .Z(
        u4_sll_454_ML_int_4__48_) );
  MUX2_X2 u4_sll_454_M1_3_49 ( .A(u4_sll_454_ML_int_3__49_), .B(
        u4_sll_454_ML_int_3__41_), .S(u4_sll_454_n19), .Z(
        u4_sll_454_ML_int_4__49_) );
  MUX2_X2 u4_sll_454_M1_3_50 ( .A(u4_sll_454_ML_int_3__50_), .B(
        u4_sll_454_ML_int_3__42_), .S(u4_sll_454_n19), .Z(
        u4_sll_454_ML_int_4__50_) );
  MUX2_X2 u4_sll_454_M1_3_51 ( .A(u4_sll_454_ML_int_3__51_), .B(
        u4_sll_454_ML_int_3__43_), .S(u4_sll_454_n19), .Z(
        u4_sll_454_ML_int_4__51_) );
  MUX2_X2 u4_sll_454_M1_3_52 ( .A(u4_sll_454_ML_int_3__52_), .B(
        u4_sll_454_ML_int_3__44_), .S(u4_sll_454_n20), .Z(
        u4_sll_454_ML_int_4__52_) );
  MUX2_X2 u4_sll_454_M1_3_53 ( .A(u4_sll_454_ML_int_3__53_), .B(
        u4_sll_454_ML_int_3__45_), .S(u4_sll_454_n20), .Z(
        u4_sll_454_ML_int_4__53_) );
  MUX2_X2 u4_sll_454_M1_3_54 ( .A(u4_sll_454_ML_int_3__54_), .B(
        u4_sll_454_ML_int_3__46_), .S(u4_sll_454_n20), .Z(
        u4_sll_454_ML_int_4__54_) );
  MUX2_X2 u4_sll_454_M1_3_55 ( .A(u4_sll_454_ML_int_3__55_), .B(
        u4_sll_454_ML_int_3__47_), .S(u4_sll_454_n20), .Z(
        u4_sll_454_ML_int_4__55_) );
  MUX2_X2 u4_sll_454_M1_3_56 ( .A(u4_sll_454_ML_int_3__56_), .B(
        u4_sll_454_ML_int_3__48_), .S(u4_sll_454_n20), .Z(
        u4_sll_454_ML_int_4__56_) );
  MUX2_X2 u4_sll_454_M1_3_57 ( .A(u4_sll_454_ML_int_3__57_), .B(
        u4_sll_454_ML_int_3__49_), .S(u4_sll_454_n20), .Z(
        u4_sll_454_ML_int_4__57_) );
  MUX2_X2 u4_sll_454_M1_3_58 ( .A(u4_sll_454_ML_int_3__58_), .B(
        u4_sll_454_ML_int_3__50_), .S(u4_sll_454_n19), .Z(
        u4_sll_454_ML_int_4__58_) );
  MUX2_X2 u4_sll_454_M1_3_59 ( .A(u4_sll_454_ML_int_3__59_), .B(
        u4_sll_454_ML_int_3__51_), .S(u4_sll_454_n19), .Z(
        u4_sll_454_ML_int_4__59_) );
  MUX2_X2 u4_sll_454_M1_3_60 ( .A(u4_sll_454_ML_int_3__60_), .B(
        u4_sll_454_ML_int_3__52_), .S(u4_sll_454_n19), .Z(
        u4_sll_454_ML_int_4__60_) );
  MUX2_X2 u4_sll_454_M1_3_61 ( .A(u4_sll_454_ML_int_3__61_), .B(
        u4_sll_454_ML_int_3__53_), .S(u4_sll_454_n19), .Z(
        u4_sll_454_ML_int_4__61_) );
  MUX2_X2 u4_sll_454_M1_3_62 ( .A(u4_sll_454_ML_int_3__62_), .B(
        u4_sll_454_ML_int_3__54_), .S(u4_sll_454_n19), .Z(
        u4_sll_454_ML_int_4__62_) );
  MUX2_X2 u4_sll_454_M1_3_63 ( .A(u4_sll_454_ML_int_3__63_), .B(
        u4_sll_454_ML_int_3__55_), .S(u4_sll_454_n20), .Z(
        u4_sll_454_ML_int_4__63_) );
  MUX2_X2 u4_sll_454_M1_3_64 ( .A(u4_sll_454_ML_int_3__64_), .B(
        u4_sll_454_ML_int_3__56_), .S(u4_sll_454_n20), .Z(
        u4_sll_454_ML_int_4__64_) );
  MUX2_X2 u4_sll_454_M1_3_65 ( .A(u4_sll_454_ML_int_3__65_), .B(
        u4_sll_454_ML_int_3__57_), .S(u4_sll_454_n20), .Z(
        u4_sll_454_ML_int_4__65_) );
  MUX2_X2 u4_sll_454_M1_3_66 ( .A(u4_sll_454_ML_int_3__66_), .B(
        u4_sll_454_ML_int_3__58_), .S(u4_sll_454_n20), .Z(
        u4_sll_454_ML_int_4__66_) );
  MUX2_X2 u4_sll_454_M1_3_67 ( .A(u4_sll_454_ML_int_3__67_), .B(
        u4_sll_454_ML_int_3__59_), .S(u4_sll_454_n20), .Z(
        u4_sll_454_ML_int_4__67_) );
  MUX2_X2 u4_sll_454_M1_3_68 ( .A(u4_sll_454_ML_int_3__68_), .B(
        u4_sll_454_ML_int_3__60_), .S(u4_sll_454_n20), .Z(
        u4_sll_454_ML_int_4__68_) );
  MUX2_X2 u4_sll_454_M1_3_69 ( .A(u4_sll_454_ML_int_3__69_), .B(
        u4_sll_454_ML_int_3__61_), .S(u4_sll_454_n20), .Z(
        u4_sll_454_ML_int_4__69_) );
  MUX2_X2 u4_sll_454_M1_3_70 ( .A(u4_sll_454_ML_int_3__70_), .B(
        u4_sll_454_ML_int_3__62_), .S(u4_sll_454_n20), .Z(
        u4_sll_454_ML_int_4__70_) );
  MUX2_X2 u4_sll_454_M1_3_71 ( .A(u4_sll_454_ML_int_3__71_), .B(
        u4_sll_454_ML_int_3__63_), .S(u4_sll_454_n20), .Z(
        u4_sll_454_ML_int_4__71_) );
  MUX2_X2 u4_sll_454_M1_3_72 ( .A(u4_sll_454_ML_int_3__72_), .B(
        u4_sll_454_ML_int_3__64_), .S(u4_sll_454_n20), .Z(
        u4_sll_454_ML_int_4__72_) );
  MUX2_X2 u4_sll_454_M1_3_73 ( .A(u4_sll_454_ML_int_3__73_), .B(
        u4_sll_454_ML_int_3__65_), .S(u4_sll_454_n20), .Z(
        u4_sll_454_ML_int_4__73_) );
  MUX2_X2 u4_sll_454_M1_3_74 ( .A(u4_sll_454_ML_int_3__74_), .B(
        u4_sll_454_ML_int_3__66_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__74_) );
  MUX2_X2 u4_sll_454_M1_3_75 ( .A(u4_sll_454_ML_int_3__75_), .B(
        u4_sll_454_ML_int_3__67_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__75_) );
  MUX2_X2 u4_sll_454_M1_3_76 ( .A(u4_sll_454_ML_int_3__76_), .B(
        u4_sll_454_ML_int_3__68_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__76_) );
  MUX2_X2 u4_sll_454_M1_3_77 ( .A(u4_sll_454_ML_int_3__77_), .B(
        u4_sll_454_ML_int_3__69_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__77_) );
  MUX2_X2 u4_sll_454_M1_3_78 ( .A(u4_sll_454_ML_int_3__78_), .B(
        u4_sll_454_ML_int_3__70_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__78_) );
  MUX2_X2 u4_sll_454_M1_3_79 ( .A(u4_sll_454_ML_int_3__79_), .B(
        u4_sll_454_ML_int_3__71_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__79_) );
  MUX2_X2 u4_sll_454_M1_3_80 ( .A(u4_sll_454_ML_int_3__80_), .B(
        u4_sll_454_ML_int_3__72_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__80_) );
  MUX2_X2 u4_sll_454_M1_3_81 ( .A(u4_sll_454_ML_int_3__81_), .B(
        u4_sll_454_ML_int_3__73_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__81_) );
  MUX2_X2 u4_sll_454_M1_3_82 ( .A(u4_sll_454_ML_int_3__82_), .B(
        u4_sll_454_ML_int_3__74_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__82_) );
  MUX2_X2 u4_sll_454_M1_3_83 ( .A(u4_sll_454_ML_int_3__83_), .B(
        u4_sll_454_ML_int_3__75_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__83_) );
  MUX2_X2 u4_sll_454_M1_3_84 ( .A(u4_sll_454_ML_int_3__84_), .B(
        u4_sll_454_ML_int_3__76_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__84_) );
  MUX2_X2 u4_sll_454_M1_3_85 ( .A(u4_sll_454_ML_int_3__85_), .B(
        u4_sll_454_ML_int_3__77_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__85_) );
  MUX2_X2 u4_sll_454_M1_3_86 ( .A(u4_sll_454_ML_int_3__86_), .B(
        u4_sll_454_ML_int_3__78_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__86_) );
  MUX2_X2 u4_sll_454_M1_3_87 ( .A(u4_sll_454_ML_int_3__87_), .B(
        u4_sll_454_ML_int_3__79_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__87_) );
  MUX2_X2 u4_sll_454_M1_3_88 ( .A(u4_sll_454_ML_int_3__88_), .B(
        u4_sll_454_ML_int_3__80_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__88_) );
  MUX2_X2 u4_sll_454_M1_3_89 ( .A(u4_sll_454_ML_int_3__89_), .B(
        u4_sll_454_ML_int_3__81_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__89_) );
  MUX2_X2 u4_sll_454_M1_3_90 ( .A(u4_sll_454_ML_int_3__90_), .B(
        u4_sll_454_ML_int_3__82_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__90_) );
  MUX2_X2 u4_sll_454_M1_3_91 ( .A(u4_sll_454_ML_int_3__91_), .B(
        u4_sll_454_ML_int_3__83_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__91_) );
  MUX2_X2 u4_sll_454_M1_3_92 ( .A(u4_sll_454_ML_int_3__92_), .B(
        u4_sll_454_ML_int_3__84_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__92_) );
  MUX2_X2 u4_sll_454_M1_3_93 ( .A(u4_sll_454_ML_int_3__93_), .B(
        u4_sll_454_ML_int_3__85_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__93_) );
  MUX2_X2 u4_sll_454_M1_3_94 ( .A(u4_sll_454_ML_int_3__94_), .B(
        u4_sll_454_ML_int_3__86_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__94_) );
  MUX2_X2 u4_sll_454_M1_3_95 ( .A(u4_sll_454_ML_int_3__95_), .B(
        u4_sll_454_ML_int_3__87_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__95_) );
  MUX2_X2 u4_sll_454_M1_3_96 ( .A(u4_sll_454_ML_int_3__96_), .B(
        u4_sll_454_ML_int_3__88_), .S(u4_sll_454_n19), .Z(
        u4_sll_454_ML_int_4__96_) );
  MUX2_X2 u4_sll_454_M1_3_97 ( .A(u4_sll_454_ML_int_3__97_), .B(
        u4_sll_454_ML_int_3__89_), .S(u4_sll_454_n19), .Z(
        u4_sll_454_ML_int_4__97_) );
  MUX2_X2 u4_sll_454_M1_3_98 ( .A(u4_sll_454_ML_int_3__98_), .B(
        u4_sll_454_ML_int_3__90_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__98_) );
  MUX2_X2 u4_sll_454_M1_3_99 ( .A(u4_sll_454_ML_int_3__99_), .B(
        u4_sll_454_ML_int_3__91_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__99_) );
  MUX2_X2 u4_sll_454_M1_3_100 ( .A(u4_sll_454_ML_int_3__100_), .B(
        u4_sll_454_ML_int_3__92_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__100_) );
  MUX2_X2 u4_sll_454_M1_3_101 ( .A(u4_sll_454_ML_int_3__101_), .B(
        u4_sll_454_ML_int_3__93_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__101_) );
  MUX2_X2 u4_sll_454_M1_3_102 ( .A(u4_sll_454_ML_int_3__102_), .B(
        u4_sll_454_ML_int_3__94_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__102_) );
  MUX2_X2 u4_sll_454_M1_3_103 ( .A(u4_sll_454_ML_int_3__103_), .B(
        u4_sll_454_ML_int_3__95_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__103_) );
  MUX2_X2 u4_sll_454_M1_3_104 ( .A(u4_sll_454_ML_int_3__104_), .B(
        u4_sll_454_ML_int_3__96_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__104_) );
  MUX2_X2 u4_sll_454_M1_3_105 ( .A(u4_sll_454_ML_int_3__105_), .B(
        u4_sll_454_ML_int_3__97_), .S(u4_sll_454_n18), .Z(
        u4_sll_454_ML_int_4__105_) );
  MUX2_X2 u4_sll_454_M1_4_16 ( .A(u4_sll_454_ML_int_4__16_), .B(
        u4_sll_454_ML_int_4__0_), .S(u4_sll_454_n32), .Z(
        u4_sll_454_ML_int_5__16_) );
  MUX2_X2 u4_sll_454_M1_4_17 ( .A(u4_sll_454_ML_int_4__17_), .B(
        u4_sll_454_ML_int_4__1_), .S(u4_sll_454_n32), .Z(
        u4_sll_454_ML_int_5__17_) );
  MUX2_X2 u4_sll_454_M1_4_18 ( .A(u4_sll_454_ML_int_4__18_), .B(
        u4_sll_454_ML_int_4__2_), .S(u4_sll_454_n31), .Z(
        u4_sll_454_ML_int_5__18_) );
  MUX2_X2 u4_sll_454_M1_4_19 ( .A(u4_sll_454_ML_int_4__19_), .B(
        u4_sll_454_ML_int_4__3_), .S(u4_sll_454_n31), .Z(
        u4_sll_454_ML_int_5__19_) );
  MUX2_X2 u4_sll_454_M1_4_20 ( .A(u4_sll_454_ML_int_4__20_), .B(
        u4_sll_454_ML_int_4__4_), .S(u4_sll_454_n31), .Z(
        u4_sll_454_ML_int_5__20_) );
  MUX2_X2 u4_sll_454_M1_4_21 ( .A(u4_sll_454_ML_int_4__21_), .B(
        u4_sll_454_ML_int_4__5_), .S(u4_sll_454_n31), .Z(
        u4_sll_454_ML_int_5__21_) );
  MUX2_X2 u4_sll_454_M1_4_22 ( .A(u4_sll_454_ML_int_4__22_), .B(
        u4_sll_454_ML_int_4__6_), .S(u4_sll_454_n31), .Z(
        u4_sll_454_ML_int_5__22_) );
  MUX2_X2 u4_sll_454_M1_4_23 ( .A(u4_sll_454_ML_int_4__23_), .B(
        u4_sll_454_ML_int_4__7_), .S(u4_sll_454_n31), .Z(
        u4_sll_454_ML_int_5__23_) );
  MUX2_X2 u4_sll_454_M1_4_24 ( .A(u4_sll_454_ML_int_4__24_), .B(
        u4_sll_454_ML_int_4__8_), .S(u4_sll_454_n31), .Z(
        u4_sll_454_ML_int_5__24_) );
  MUX2_X2 u4_sll_454_M1_4_25 ( .A(u4_sll_454_ML_int_4__25_), .B(
        u4_sll_454_ML_int_4__9_), .S(u4_sll_454_n31), .Z(
        u4_sll_454_ML_int_5__25_) );
  MUX2_X2 u4_sll_454_M1_4_26 ( .A(u4_sll_454_ML_int_4__26_), .B(
        u4_sll_454_ML_int_4__10_), .S(u4_sll_454_n31), .Z(
        u4_sll_454_ML_int_5__26_) );
  MUX2_X2 u4_sll_454_M1_4_27 ( .A(u4_sll_454_ML_int_4__27_), .B(
        u4_sll_454_ML_int_4__11_), .S(u4_sll_454_n32), .Z(
        u4_sll_454_ML_int_5__27_) );
  MUX2_X2 u4_sll_454_M1_4_28 ( .A(u4_sll_454_ML_int_4__28_), .B(
        u4_sll_454_ML_int_4__12_), .S(u4_sll_454_n32), .Z(
        u4_sll_454_ML_int_5__28_) );
  MUX2_X2 u4_sll_454_M1_4_29 ( .A(u4_sll_454_ML_int_4__29_), .B(
        u4_sll_454_ML_int_4__13_), .S(u4_sll_454_n32), .Z(
        u4_sll_454_ML_int_5__29_) );
  MUX2_X2 u4_sll_454_M1_4_30 ( .A(u4_sll_454_ML_int_4__30_), .B(
        u4_sll_454_ML_int_4__14_), .S(u4_sll_454_n32), .Z(
        u4_sll_454_ML_int_5__30_) );
  MUX2_X2 u4_sll_454_M1_4_31 ( .A(u4_sll_454_ML_int_4__31_), .B(
        u4_sll_454_ML_int_4__15_), .S(u4_sll_454_n32), .Z(
        u4_sll_454_ML_int_5__31_) );
  MUX2_X2 u4_sll_454_M1_4_32 ( .A(u4_sll_454_ML_int_4__32_), .B(
        u4_sll_454_ML_int_4__16_), .S(u4_sll_454_n32), .Z(
        u4_sll_454_ML_int_5__32_) );
  MUX2_X2 u4_sll_454_M1_4_33 ( .A(u4_sll_454_ML_int_4__33_), .B(
        u4_sll_454_ML_int_4__17_), .S(u4_sll_454_n32), .Z(
        u4_sll_454_ML_int_5__33_) );
  MUX2_X2 u4_sll_454_M1_4_34 ( .A(u4_sll_454_ML_int_4__34_), .B(
        u4_sll_454_ML_int_4__18_), .S(u4_sll_454_n32), .Z(
        u4_sll_454_ML_int_5__34_) );
  MUX2_X2 u4_sll_454_M1_4_35 ( .A(u4_sll_454_ML_int_4__35_), .B(
        u4_sll_454_ML_int_4__19_), .S(u4_sll_454_n32), .Z(
        u4_sll_454_ML_int_5__35_) );
  MUX2_X2 u4_sll_454_M1_4_36 ( .A(u4_sll_454_ML_int_4__36_), .B(
        u4_sll_454_ML_int_4__20_), .S(u4_sll_454_n32), .Z(
        u4_sll_454_ML_int_5__36_) );
  MUX2_X2 u4_sll_454_M1_4_37 ( .A(u4_sll_454_ML_int_4__37_), .B(
        u4_sll_454_ML_int_4__21_), .S(u4_sll_454_n32), .Z(
        u4_sll_454_ML_int_5__37_) );
  MUX2_X2 u4_sll_454_M1_4_38 ( .A(u4_sll_454_ML_int_4__38_), .B(
        u4_sll_454_ML_int_4__22_), .S(u4_sll_454_n28), .Z(
        u4_sll_454_ML_int_5__38_) );
  MUX2_X2 u4_sll_454_M1_4_39 ( .A(u4_sll_454_ML_int_4__39_), .B(
        u4_sll_454_ML_int_4__23_), .S(u4_sll_454_n27), .Z(
        u4_sll_454_ML_int_5__39_) );
  MUX2_X2 u4_sll_454_M1_4_40 ( .A(u4_sll_454_ML_int_4__40_), .B(
        u4_sll_454_ML_int_4__24_), .S(u4_sll_454_n27), .Z(
        u4_sll_454_ML_int_5__40_) );
  MUX2_X2 u4_sll_454_M1_4_41 ( .A(u4_sll_454_ML_int_4__41_), .B(
        u4_sll_454_ML_int_4__25_), .S(u4_sll_454_n27), .Z(
        u4_sll_454_ML_int_5__41_) );
  MUX2_X2 u4_sll_454_M1_4_42 ( .A(u4_sll_454_ML_int_4__42_), .B(
        u4_sll_454_ML_int_4__26_), .S(u4_sll_454_n27), .Z(
        u4_sll_454_ML_int_5__42_) );
  MUX2_X2 u4_sll_454_M1_4_43 ( .A(u4_sll_454_ML_int_4__43_), .B(
        u4_sll_454_ML_int_4__27_), .S(u4_sll_454_n27), .Z(
        u4_sll_454_ML_int_5__43_) );
  MUX2_X2 u4_sll_454_M1_4_44 ( .A(u4_sll_454_ML_int_4__44_), .B(
        u4_sll_454_ML_int_4__28_), .S(u4_sll_454_n32), .Z(
        u4_sll_454_ML_int_5__44_) );
  MUX2_X2 u4_sll_454_M1_4_45 ( .A(u4_sll_454_ML_int_4__45_), .B(
        u4_sll_454_ML_int_4__29_), .S(u4_sll_454_n32), .Z(
        u4_sll_454_ML_int_5__45_) );
  MUX2_X2 u4_sll_454_M1_4_46 ( .A(u4_sll_454_ML_int_4__46_), .B(
        u4_sll_454_ML_int_4__30_), .S(u4_sll_454_n32), .Z(
        u4_sll_454_ML_int_5__46_) );
  MUX2_X2 u4_sll_454_M1_4_47 ( .A(u4_sll_454_ML_int_4__47_), .B(
        u4_sll_454_ML_int_4__31_), .S(u4_sll_454_n32), .Z(
        u4_sll_454_ML_int_5__47_) );
  MUX2_X2 u4_sll_454_M1_4_48 ( .A(u4_sll_454_ML_int_4__48_), .B(
        u4_sll_454_ML_int_4__32_), .S(u4_sll_454_n32), .Z(
        u4_sll_454_ML_int_5__48_) );
  MUX2_X2 u4_sll_454_M1_4_49 ( .A(u4_sll_454_ML_int_4__49_), .B(
        u4_sll_454_ML_int_4__33_), .S(u4_sll_454_n30), .Z(
        u4_sll_454_ML_int_5__49_) );
  MUX2_X2 u4_sll_454_M1_4_50 ( .A(u4_sll_454_ML_int_4__50_), .B(
        u4_sll_454_ML_int_4__34_), .S(u4_sll_454_n30), .Z(
        u4_sll_454_ML_int_5__50_) );
  MUX2_X2 u4_sll_454_M1_4_51 ( .A(u4_sll_454_ML_int_4__51_), .B(
        u4_sll_454_ML_int_4__35_), .S(u4_sll_454_n30), .Z(
        u4_sll_454_ML_int_5__51_) );
  MUX2_X2 u4_sll_454_M1_4_52 ( .A(u4_sll_454_ML_int_4__52_), .B(
        u4_sll_454_ML_int_4__36_), .S(u4_sll_454_n30), .Z(
        u4_sll_454_ML_int_5__52_) );
  MUX2_X2 u4_sll_454_M1_4_53 ( .A(u4_sll_454_ML_int_4__53_), .B(
        u4_sll_454_ML_int_4__37_), .S(u4_sll_454_n30), .Z(
        u4_sll_454_ML_int_5__53_) );
  MUX2_X2 u4_sll_454_M1_4_54 ( .A(u4_sll_454_ML_int_4__54_), .B(
        u4_sll_454_ML_int_4__38_), .S(u4_sll_454_n29), .Z(
        u4_sll_454_ML_int_5__54_) );
  MUX2_X2 u4_sll_454_M1_4_55 ( .A(u4_sll_454_ML_int_4__55_), .B(
        u4_sll_454_ML_int_4__39_), .S(u4_sll_454_n29), .Z(
        u4_sll_454_ML_int_5__55_) );
  MUX2_X2 u4_sll_454_M1_4_56 ( .A(u4_sll_454_ML_int_4__56_), .B(
        u4_sll_454_ML_int_4__40_), .S(u4_sll_454_n29), .Z(
        u4_sll_454_ML_int_5__56_) );
  MUX2_X2 u4_sll_454_M1_4_57 ( .A(u4_sll_454_ML_int_4__57_), .B(
        u4_sll_454_ML_int_4__41_), .S(u4_sll_454_n29), .Z(
        u4_sll_454_ML_int_5__57_) );
  MUX2_X2 u4_sll_454_M1_4_58 ( .A(u4_sll_454_ML_int_4__58_), .B(
        u4_sll_454_ML_int_4__42_), .S(u4_sll_454_n29), .Z(
        u4_sll_454_ML_int_5__58_) );
  MUX2_X2 u4_sll_454_M1_4_59 ( .A(u4_sll_454_ML_int_4__59_), .B(
        u4_sll_454_ML_int_4__43_), .S(u4_sll_454_n29), .Z(
        u4_sll_454_ML_int_5__59_) );
  MUX2_X2 u4_sll_454_M1_4_60 ( .A(u4_sll_454_ML_int_4__60_), .B(
        u4_sll_454_ML_int_4__44_), .S(u4_sll_454_n30), .Z(
        u4_sll_454_ML_int_5__60_) );
  MUX2_X2 u4_sll_454_M1_4_61 ( .A(u4_sll_454_ML_int_4__61_), .B(
        u4_sll_454_ML_int_4__45_), .S(u4_sll_454_n30), .Z(
        u4_sll_454_ML_int_5__61_) );
  MUX2_X2 u4_sll_454_M1_4_62 ( .A(u4_sll_454_ML_int_4__62_), .B(
        u4_sll_454_ML_int_4__46_), .S(u4_sll_454_n30), .Z(
        u4_sll_454_ML_int_5__62_) );
  MUX2_X2 u4_sll_454_M1_4_63 ( .A(u4_sll_454_ML_int_4__63_), .B(
        u4_sll_454_ML_int_4__47_), .S(u4_sll_454_n30), .Z(
        u4_sll_454_ML_int_5__63_) );
  MUX2_X2 u4_sll_454_M1_4_64 ( .A(u4_sll_454_ML_int_4__64_), .B(
        u4_sll_454_ML_int_4__48_), .S(u4_sll_454_n30), .Z(
        u4_sll_454_ML_int_5__64_) );
  MUX2_X2 u4_sll_454_M1_4_65 ( .A(u4_sll_454_ML_int_4__65_), .B(
        u4_sll_454_ML_int_4__49_), .S(u4_sll_454_n30), .Z(
        u4_sll_454_ML_int_5__65_) );
  MUX2_X2 u4_sll_454_M1_4_66 ( .A(u4_sll_454_ML_int_4__66_), .B(
        u4_sll_454_ML_int_4__50_), .S(u4_sll_454_n30), .Z(
        u4_sll_454_ML_int_5__66_) );
  MUX2_X2 u4_sll_454_M1_4_67 ( .A(u4_sll_454_ML_int_4__67_), .B(
        u4_sll_454_ML_int_4__51_), .S(u4_sll_454_n30), .Z(
        u4_sll_454_ML_int_5__67_) );
  MUX2_X2 u4_sll_454_M1_4_68 ( .A(u4_sll_454_ML_int_4__68_), .B(
        u4_sll_454_ML_int_4__52_), .S(u4_sll_454_n30), .Z(
        u4_sll_454_ML_int_5__68_) );
  MUX2_X2 u4_sll_454_M1_4_69 ( .A(u4_sll_454_ML_int_4__69_), .B(
        u4_sll_454_ML_int_4__53_), .S(u4_sll_454_n30), .Z(
        u4_sll_454_ML_int_5__69_) );
  MUX2_X2 u4_sll_454_M1_4_70 ( .A(u4_sll_454_ML_int_4__70_), .B(
        u4_sll_454_ML_int_4__54_), .S(u4_sll_454_n30), .Z(
        u4_sll_454_ML_int_5__70_) );
  MUX2_X2 u4_sll_454_M1_4_71 ( .A(u4_sll_454_ML_int_4__71_), .B(
        u4_sll_454_ML_int_4__55_), .S(u4_sll_454_n31), .Z(
        u4_sll_454_ML_int_5__71_) );
  MUX2_X2 u4_sll_454_M1_4_72 ( .A(u4_sll_454_ML_int_4__72_), .B(
        u4_sll_454_ML_int_4__56_), .S(u4_sll_454_n31), .Z(
        u4_sll_454_ML_int_5__72_) );
  MUX2_X2 u4_sll_454_M1_4_73 ( .A(u4_sll_454_ML_int_4__73_), .B(
        u4_sll_454_ML_int_4__57_), .S(u4_sll_454_n31), .Z(
        u4_sll_454_ML_int_5__73_) );
  MUX2_X2 u4_sll_454_M1_4_74 ( .A(u4_sll_454_ML_int_4__74_), .B(
        u4_sll_454_ML_int_4__58_), .S(u4_sll_454_n31), .Z(
        u4_sll_454_ML_int_5__74_) );
  MUX2_X2 u4_sll_454_M1_4_75 ( .A(u4_sll_454_ML_int_4__75_), .B(
        u4_sll_454_ML_int_4__59_), .S(u4_sll_454_n31), .Z(
        u4_sll_454_ML_int_5__75_) );
  MUX2_X2 u4_sll_454_M1_4_76 ( .A(u4_sll_454_ML_int_4__76_), .B(
        u4_sll_454_ML_int_4__60_), .S(u4_sll_454_n31), .Z(
        u4_sll_454_ML_int_5__76_) );
  MUX2_X2 u4_sll_454_M1_4_77 ( .A(u4_sll_454_ML_int_4__77_), .B(
        u4_sll_454_ML_int_4__61_), .S(u4_sll_454_n31), .Z(
        u4_sll_454_ML_int_5__77_) );
  MUX2_X2 u4_sll_454_M1_4_78 ( .A(u4_sll_454_ML_int_4__78_), .B(
        u4_sll_454_ML_int_4__62_), .S(u4_sll_454_n31), .Z(
        u4_sll_454_ML_int_5__78_) );
  MUX2_X2 u4_sll_454_M1_4_79 ( .A(u4_sll_454_ML_int_4__79_), .B(
        u4_sll_454_ML_int_4__63_), .S(u4_sll_454_n31), .Z(
        u4_sll_454_ML_int_5__79_) );
  MUX2_X2 u4_sll_454_M1_4_80 ( .A(u4_sll_454_ML_int_4__80_), .B(
        u4_sll_454_ML_int_4__64_), .S(u4_sll_454_n30), .Z(
        u4_sll_454_ML_int_5__80_) );
  MUX2_X2 u4_sll_454_M1_4_81 ( .A(u4_sll_454_ML_int_4__81_), .B(
        u4_sll_454_ML_int_4__65_), .S(u4_sll_454_n30), .Z(
        u4_sll_454_ML_int_5__81_) );
  MUX2_X2 u4_sll_454_M1_4_82 ( .A(u4_sll_454_ML_int_4__82_), .B(
        u4_sll_454_ML_int_4__66_), .S(u4_sll_454_n27), .Z(
        u4_sll_454_ML_int_5__82_) );
  MUX2_X2 u4_sll_454_M1_4_83 ( .A(u4_sll_454_ML_int_4__83_), .B(
        u4_sll_454_ML_int_4__67_), .S(u4_sll_454_n27), .Z(
        u4_sll_454_ML_int_5__83_) );
  MUX2_X2 u4_sll_454_M1_4_84 ( .A(u4_sll_454_ML_int_4__84_), .B(
        u4_sll_454_ML_int_4__68_), .S(u4_sll_454_n27), .Z(
        u4_sll_454_ML_int_5__84_) );
  MUX2_X2 u4_sll_454_M1_4_85 ( .A(u4_sll_454_ML_int_4__85_), .B(
        u4_sll_454_ML_int_4__69_), .S(u4_sll_454_n27), .Z(
        u4_sll_454_ML_int_5__85_) );
  MUX2_X2 u4_sll_454_M1_4_86 ( .A(u4_sll_454_ML_int_4__86_), .B(
        u4_sll_454_ML_int_4__70_), .S(u4_sll_454_n27), .Z(
        u4_sll_454_ML_int_5__86_) );
  MUX2_X2 u4_sll_454_M1_4_87 ( .A(u4_sll_454_ML_int_4__87_), .B(
        u4_sll_454_ML_int_4__71_), .S(u4_sll_454_n27), .Z(
        u4_sll_454_ML_int_5__87_) );
  MUX2_X2 u4_sll_454_M1_4_88 ( .A(u4_sll_454_ML_int_4__88_), .B(
        u4_sll_454_ML_int_4__72_), .S(u4_sll_454_n27), .Z(
        u4_sll_454_ML_int_5__88_) );
  MUX2_X2 u4_sll_454_M1_4_89 ( .A(u4_sll_454_ML_int_4__89_), .B(
        u4_sll_454_ML_int_4__73_), .S(u4_sll_454_n28), .Z(
        u4_sll_454_ML_int_5__89_) );
  MUX2_X2 u4_sll_454_M1_4_90 ( .A(u4_sll_454_ML_int_4__90_), .B(
        u4_sll_454_ML_int_4__74_), .S(u4_sll_454_n27), .Z(
        u4_sll_454_ML_int_5__90_) );
  MUX2_X2 u4_sll_454_M1_4_91 ( .A(u4_sll_454_ML_int_4__91_), .B(
        u4_sll_454_ML_int_4__75_), .S(u4_sll_454_n28), .Z(
        u4_sll_454_ML_int_5__91_) );
  MUX2_X2 u4_sll_454_M1_4_92 ( .A(u4_sll_454_ML_int_4__92_), .B(
        u4_sll_454_ML_int_4__76_), .S(u4_sll_454_n27), .Z(
        u4_sll_454_ML_int_5__92_) );
  MUX2_X2 u4_sll_454_M1_4_93 ( .A(u4_sll_454_ML_int_4__93_), .B(
        u4_sll_454_ML_int_4__77_), .S(u4_sll_454_n29), .Z(
        u4_sll_454_ML_int_5__93_) );
  MUX2_X2 u4_sll_454_M1_4_94 ( .A(u4_sll_454_ML_int_4__94_), .B(
        u4_sll_454_ML_int_4__78_), .S(u4_sll_454_n29), .Z(
        u4_sll_454_ML_int_5__94_) );
  MUX2_X2 u4_sll_454_M1_4_95 ( .A(u4_sll_454_ML_int_4__95_), .B(
        u4_sll_454_ML_int_4__79_), .S(u4_sll_454_n29), .Z(
        u4_sll_454_ML_int_5__95_) );
  MUX2_X2 u4_sll_454_M1_4_96 ( .A(u4_sll_454_ML_int_4__96_), .B(
        u4_sll_454_ML_int_4__80_), .S(u4_sll_454_n29), .Z(
        u4_sll_454_ML_int_5__96_) );
  MUX2_X2 u4_sll_454_M1_4_97 ( .A(u4_sll_454_ML_int_4__97_), .B(
        u4_sll_454_ML_int_4__81_), .S(u4_sll_454_n29), .Z(
        u4_sll_454_ML_int_5__97_) );
  MUX2_X2 u4_sll_454_M1_4_98 ( .A(u4_sll_454_ML_int_4__98_), .B(
        u4_sll_454_ML_int_4__82_), .S(u4_sll_454_n29), .Z(
        u4_sll_454_ML_int_5__98_) );
  MUX2_X2 u4_sll_454_M1_4_99 ( .A(u4_sll_454_ML_int_4__99_), .B(
        u4_sll_454_ML_int_4__83_), .S(u4_sll_454_n29), .Z(
        u4_sll_454_ML_int_5__99_) );
  MUX2_X2 u4_sll_454_M1_4_100 ( .A(u4_sll_454_ML_int_4__100_), .B(
        u4_sll_454_ML_int_4__84_), .S(u4_sll_454_n29), .Z(
        u4_sll_454_ML_int_5__100_) );
  MUX2_X2 u4_sll_454_M1_4_101 ( .A(u4_sll_454_ML_int_4__101_), .B(
        u4_sll_454_ML_int_4__85_), .S(u4_sll_454_n29), .Z(
        u4_sll_454_ML_int_5__101_) );
  MUX2_X2 u4_sll_454_M1_4_102 ( .A(u4_sll_454_ML_int_4__102_), .B(
        u4_sll_454_ML_int_4__86_), .S(u4_sll_454_n29), .Z(
        u4_sll_454_ML_int_5__102_) );
  MUX2_X2 u4_sll_454_M1_4_103 ( .A(u4_sll_454_ML_int_4__103_), .B(
        u4_sll_454_ML_int_4__87_), .S(u4_sll_454_n28), .Z(
        u4_sll_454_ML_int_5__103_) );
  MUX2_X2 u4_sll_454_M1_4_104 ( .A(u4_sll_454_ML_int_4__104_), .B(
        u4_sll_454_ML_int_4__88_), .S(u4_sll_454_n29), .Z(
        u4_sll_454_ML_int_5__104_) );
  MUX2_X2 u4_sll_454_M1_4_105 ( .A(u4_sll_454_ML_int_4__105_), .B(
        u4_sll_454_ML_int_4__89_), .S(u4_sll_454_n29), .Z(
        u4_sll_454_ML_int_5__105_) );
  MUX2_X2 u4_sll_454_M1_5_32 ( .A(u4_sll_454_ML_int_5__32_), .B(
        u4_sll_454_ML_int_5__0_), .S(u4_sll_454_n44), .Z(
        u4_sll_454_ML_int_6__32_) );
  MUX2_X2 u4_sll_454_M1_5_33 ( .A(u4_sll_454_ML_int_5__33_), .B(
        u4_sll_454_ML_int_5__1_), .S(u4_sll_454_n44), .Z(
        u4_sll_454_ML_int_6__33_) );
  MUX2_X2 u4_sll_454_M1_5_34 ( .A(u4_sll_454_ML_int_5__34_), .B(
        u4_sll_454_ML_int_5__2_), .S(u4_sll_454_n44), .Z(
        u4_sll_454_ML_int_6__34_) );
  MUX2_X2 u4_sll_454_M1_5_35 ( .A(u4_sll_454_ML_int_5__35_), .B(
        u4_sll_454_ML_int_5__3_), .S(u4_sll_454_n44), .Z(
        u4_sll_454_ML_int_6__35_) );
  MUX2_X2 u4_sll_454_M1_5_36 ( .A(u4_sll_454_ML_int_5__36_), .B(
        u4_sll_454_ML_int_5__4_), .S(u4_sll_454_n44), .Z(
        u4_sll_454_ML_int_6__36_) );
  MUX2_X2 u4_sll_454_M1_5_37 ( .A(u4_sll_454_ML_int_5__37_), .B(
        u4_sll_454_ML_int_5__5_), .S(u4_sll_454_n44), .Z(
        u4_sll_454_ML_int_6__37_) );
  MUX2_X2 u4_sll_454_M1_5_38 ( .A(u4_sll_454_ML_int_5__38_), .B(
        u4_sll_454_ML_int_5__6_), .S(u4_sll_454_n45), .Z(
        u4_sll_454_ML_int_6__38_) );
  MUX2_X2 u4_sll_454_M1_5_39 ( .A(u4_sll_454_ML_int_5__39_), .B(
        u4_sll_454_ML_int_5__7_), .S(u4_sll_454_n45), .Z(
        u4_sll_454_ML_int_6__39_) );
  MUX2_X2 u4_sll_454_M1_5_40 ( .A(u4_sll_454_ML_int_5__40_), .B(
        u4_sll_454_ML_int_5__8_), .S(u4_sll_454_n45), .Z(
        u4_sll_454_ML_int_6__40_) );
  MUX2_X2 u4_sll_454_M1_5_41 ( .A(u4_sll_454_ML_int_5__41_), .B(
        u4_sll_454_ML_int_5__9_), .S(u4_sll_454_n45), .Z(
        u4_sll_454_ML_int_6__41_) );
  MUX2_X2 u4_sll_454_M1_5_42 ( .A(u4_sll_454_ML_int_5__42_), .B(
        u4_sll_454_ML_int_5__10_), .S(u4_sll_454_n45), .Z(
        u4_sll_454_ML_int_6__42_) );
  MUX2_X2 u4_sll_454_M1_5_43 ( .A(u4_sll_454_ML_int_5__43_), .B(
        u4_sll_454_ML_int_5__11_), .S(u4_sll_454_n45), .Z(
        u4_sll_454_ML_int_6__43_) );
  MUX2_X2 u4_sll_454_M1_5_44 ( .A(u4_sll_454_ML_int_5__44_), .B(
        u4_sll_454_ML_int_5__12_), .S(u4_sll_454_n45), .Z(
        u4_sll_454_ML_int_6__44_) );
  MUX2_X2 u4_sll_454_M1_5_45 ( .A(u4_sll_454_ML_int_5__45_), .B(
        u4_sll_454_ML_int_5__13_), .S(u4_sll_454_n45), .Z(
        u4_sll_454_ML_int_6__45_) );
  MUX2_X2 u4_sll_454_M1_5_46 ( .A(u4_sll_454_ML_int_5__46_), .B(
        u4_sll_454_ML_int_5__14_), .S(u4_sll_454_n45), .Z(
        u4_sll_454_ML_int_6__46_) );
  MUX2_X2 u4_sll_454_M1_5_47 ( .A(u4_sll_454_ML_int_5__47_), .B(
        u4_sll_454_ML_int_5__15_), .S(u4_sll_454_n45), .Z(
        u4_sll_454_ML_int_6__47_) );
  MUX2_X2 u4_sll_454_M1_5_48 ( .A(u4_sll_454_ML_int_5__48_), .B(
        u4_sll_454_ML_int_5__16_), .S(u4_sll_454_n45), .Z(
        u4_sll_454_ML_int_6__48_) );
  MUX2_X2 u4_sll_454_M1_5_49 ( .A(u4_sll_454_ML_int_5__49_), .B(
        u4_sll_454_ML_int_5__17_), .S(u4_sll_454_n45), .Z(
        u4_sll_454_ML_int_6__49_) );
  MUX2_X2 u4_sll_454_M1_5_50 ( .A(u4_sll_454_ML_int_5__50_), .B(
        u4_sll_454_ML_int_5__18_), .S(u4_sll_454_n45), .Z(
        u4_sll_454_ML_int_6__50_) );
  MUX2_X2 u4_sll_454_M1_5_51 ( .A(u4_sll_454_ML_int_5__51_), .B(
        u4_sll_454_ML_int_5__19_), .S(u4_sll_454_n45), .Z(
        u4_sll_454_ML_int_6__51_) );
  MUX2_X2 u4_sll_454_M1_5_52 ( .A(u4_sll_454_ML_int_5__52_), .B(
        u4_sll_454_ML_int_5__20_), .S(u4_sll_454_n45), .Z(
        u4_sll_454_ML_int_6__52_) );
  MUX2_X2 u4_sll_454_M1_5_53 ( .A(u4_sll_454_ML_int_5__53_), .B(
        u4_sll_454_ML_int_5__21_), .S(u4_sll_454_n45), .Z(
        u4_sll_454_ML_int_6__53_) );
  MUX2_X2 u4_sll_454_M1_5_54 ( .A(u4_sll_454_ML_int_5__54_), .B(
        u4_sll_454_ML_int_5__22_), .S(u4_sll_454_n45), .Z(
        u4_sll_454_ML_int_6__54_) );
  MUX2_X2 u4_sll_454_M1_5_55 ( .A(u4_sll_454_ML_int_5__55_), .B(
        u4_sll_454_ML_int_5__23_), .S(u4_sll_454_n45), .Z(
        u4_sll_454_ML_int_6__55_) );
  MUX2_X2 u4_sll_454_M1_5_56 ( .A(u4_sll_454_ML_int_5__56_), .B(
        u4_sll_454_ML_int_5__24_), .S(u4_sll_454_n46), .Z(
        u4_sll_454_ML_int_6__56_) );
  MUX2_X2 u4_sll_454_M1_5_57 ( .A(u4_sll_454_ML_int_5__57_), .B(
        u4_sll_454_ML_int_5__25_), .S(u4_sll_454_n46), .Z(
        u4_sll_454_ML_int_6__57_) );
  MUX2_X2 u4_sll_454_M1_5_58 ( .A(u4_sll_454_ML_int_5__58_), .B(
        u4_sll_454_ML_int_5__26_), .S(u4_sll_454_n46), .Z(
        u4_sll_454_ML_int_6__58_) );
  MUX2_X2 u4_sll_454_M1_5_59 ( .A(u4_sll_454_ML_int_5__59_), .B(
        u4_sll_454_ML_int_5__27_), .S(u4_sll_454_n46), .Z(
        u4_sll_454_ML_int_6__59_) );
  MUX2_X2 u4_sll_454_M1_5_60 ( .A(u4_sll_454_ML_int_5__60_), .B(
        u4_sll_454_ML_int_5__28_), .S(u4_sll_454_n46), .Z(
        u4_sll_454_ML_int_6__60_) );
  MUX2_X2 u4_sll_454_M1_5_61 ( .A(u4_sll_454_ML_int_5__61_), .B(
        u4_sll_454_ML_int_5__29_), .S(u4_sll_454_n46), .Z(
        u4_sll_454_ML_int_6__61_) );
  MUX2_X2 u4_sll_454_M1_5_62 ( .A(u4_sll_454_ML_int_5__62_), .B(
        u4_sll_454_ML_int_5__30_), .S(u4_sll_454_n46), .Z(
        u4_sll_454_ML_int_6__62_) );
  MUX2_X2 u4_sll_454_M1_5_63 ( .A(u4_sll_454_ML_int_5__63_), .B(
        u4_sll_454_ML_int_5__31_), .S(u4_sll_454_n46), .Z(
        u4_sll_454_ML_int_6__63_) );
  MUX2_X2 u4_sll_454_M1_5_64 ( .A(u4_sll_454_ML_int_5__64_), .B(
        u4_sll_454_ML_int_5__32_), .S(u4_sll_454_n46), .Z(
        u4_sll_454_ML_int_6__64_) );
  MUX2_X2 u4_sll_454_M1_5_65 ( .A(u4_sll_454_ML_int_5__65_), .B(
        u4_sll_454_ML_int_5__33_), .S(u4_sll_454_n46), .Z(
        u4_sll_454_ML_int_6__65_) );
  MUX2_X2 u4_sll_454_M1_5_66 ( .A(u4_sll_454_ML_int_5__66_), .B(
        u4_sll_454_ML_int_5__34_), .S(u4_sll_454_n46), .Z(
        u4_sll_454_ML_int_6__66_) );
  MUX2_X2 u4_sll_454_M1_5_67 ( .A(u4_sll_454_ML_int_5__67_), .B(
        u4_sll_454_ML_int_5__35_), .S(u4_sll_454_n46), .Z(
        u4_sll_454_ML_int_6__67_) );
  MUX2_X2 u4_sll_454_M1_5_68 ( .A(u4_sll_454_ML_int_5__68_), .B(
        u4_sll_454_ML_int_5__36_), .S(u4_sll_454_n46), .Z(
        u4_sll_454_ML_int_6__68_) );
  MUX2_X2 u4_sll_454_M1_5_69 ( .A(u4_sll_454_ML_int_5__69_), .B(
        u4_sll_454_ML_int_5__37_), .S(u4_sll_454_n46), .Z(
        u4_sll_454_ML_int_6__69_) );
  MUX2_X2 u4_sll_454_M1_5_70 ( .A(u4_sll_454_ML_int_5__70_), .B(
        u4_sll_454_ML_int_5__38_), .S(u4_sll_454_n46), .Z(
        u4_sll_454_ML_int_6__70_) );
  MUX2_X2 u4_sll_454_M1_5_71 ( .A(u4_sll_454_ML_int_5__71_), .B(
        u4_sll_454_ML_int_5__39_), .S(u4_sll_454_n46), .Z(
        u4_sll_454_ML_int_6__71_) );
  MUX2_X2 u4_sll_454_M1_5_72 ( .A(u4_sll_454_ML_int_5__72_), .B(
        u4_sll_454_ML_int_5__40_), .S(u4_sll_454_n46), .Z(
        u4_sll_454_ML_int_6__72_) );
  MUX2_X2 u4_sll_454_M1_5_73 ( .A(u4_sll_454_ML_int_5__73_), .B(
        u4_sll_454_ML_int_5__41_), .S(u4_sll_454_n46), .Z(
        u4_sll_454_ML_int_6__73_) );
  MUX2_X2 u4_sll_454_M1_5_74 ( .A(u4_sll_454_ML_int_5__74_), .B(
        u4_sll_454_ML_int_5__42_), .S(u4_sll_454_n47), .Z(
        u4_sll_454_ML_int_6__74_) );
  MUX2_X2 u4_sll_454_M1_5_75 ( .A(u4_sll_454_ML_int_5__75_), .B(
        u4_sll_454_ML_int_5__43_), .S(u4_sll_454_n47), .Z(
        u4_sll_454_ML_int_6__75_) );
  MUX2_X2 u4_sll_454_M1_5_76 ( .A(u4_sll_454_ML_int_5__76_), .B(
        u4_sll_454_ML_int_5__44_), .S(u4_sll_454_n47), .Z(
        u4_sll_454_ML_int_6__76_) );
  MUX2_X2 u4_sll_454_M1_5_77 ( .A(u4_sll_454_ML_int_5__77_), .B(
        u4_sll_454_ML_int_5__45_), .S(u4_sll_454_n47), .Z(
        u4_sll_454_ML_int_6__77_) );
  MUX2_X2 u4_sll_454_M1_5_78 ( .A(u4_sll_454_ML_int_5__78_), .B(
        u4_sll_454_ML_int_5__46_), .S(u4_sll_454_n47), .Z(
        u4_sll_454_ML_int_6__78_) );
  MUX2_X2 u4_sll_454_M1_5_79 ( .A(u4_sll_454_ML_int_5__79_), .B(
        u4_sll_454_ML_int_5__47_), .S(u4_sll_454_n47), .Z(
        u4_sll_454_ML_int_6__79_) );
  MUX2_X2 u4_sll_454_M1_5_80 ( .A(u4_sll_454_ML_int_5__80_), .B(
        u4_sll_454_ML_int_5__48_), .S(u4_sll_454_n47), .Z(
        u4_sll_454_ML_int_6__80_) );
  MUX2_X2 u4_sll_454_M1_5_81 ( .A(u4_sll_454_ML_int_5__81_), .B(
        u4_sll_454_ML_int_5__49_), .S(u4_sll_454_n47), .Z(
        u4_sll_454_ML_int_6__81_) );
  MUX2_X2 u4_sll_454_M1_5_82 ( .A(u4_sll_454_ML_int_5__82_), .B(
        u4_sll_454_ML_int_5__50_), .S(u4_sll_454_n47), .Z(
        u4_sll_454_ML_int_6__82_) );
  MUX2_X2 u4_sll_454_M1_5_83 ( .A(u4_sll_454_ML_int_5__83_), .B(
        u4_sll_454_ML_int_5__51_), .S(u4_sll_454_n47), .Z(
        u4_sll_454_ML_int_6__83_) );
  MUX2_X2 u4_sll_454_M1_5_84 ( .A(u4_sll_454_ML_int_5__84_), .B(
        u4_sll_454_ML_int_5__52_), .S(u4_sll_454_n47), .Z(
        u4_sll_454_ML_int_6__84_) );
  MUX2_X2 u4_sll_454_M1_5_85 ( .A(u4_sll_454_ML_int_5__85_), .B(
        u4_sll_454_ML_int_5__53_), .S(u4_sll_454_n47), .Z(
        u4_sll_454_ML_int_6__85_) );
  MUX2_X2 u4_sll_454_M1_5_86 ( .A(u4_sll_454_ML_int_5__86_), .B(
        u4_sll_454_ML_int_5__54_), .S(u4_sll_454_n47), .Z(
        u4_sll_454_ML_int_6__86_) );
  MUX2_X2 u4_sll_454_M1_5_87 ( .A(u4_sll_454_ML_int_5__87_), .B(
        u4_sll_454_ML_int_5__55_), .S(u4_sll_454_n47), .Z(
        u4_sll_454_ML_int_6__87_) );
  MUX2_X2 u4_sll_454_M1_5_88 ( .A(u4_sll_454_ML_int_5__88_), .B(
        u4_sll_454_ML_int_5__56_), .S(u4_sll_454_n47), .Z(
        u4_sll_454_ML_int_6__88_) );
  MUX2_X2 u4_sll_454_M1_5_89 ( .A(u4_sll_454_ML_int_5__89_), .B(
        u4_sll_454_ML_int_5__57_), .S(u4_sll_454_n47), .Z(
        u4_sll_454_ML_int_6__89_) );
  MUX2_X2 u4_sll_454_M1_5_90 ( .A(u4_sll_454_ML_int_5__90_), .B(
        u4_sll_454_ML_int_5__58_), .S(u4_sll_454_n47), .Z(
        u4_sll_454_ML_int_6__90_) );
  MUX2_X2 u4_sll_454_M1_5_91 ( .A(u4_sll_454_ML_int_5__91_), .B(
        u4_sll_454_ML_int_5__59_), .S(u4_sll_454_n47), .Z(
        u4_sll_454_ML_int_6__91_) );
  MUX2_X2 u4_sll_454_M1_5_92 ( .A(u4_sll_454_ML_int_5__92_), .B(
        u4_sll_454_ML_int_5__60_), .S(u4_sll_454_n43), .Z(
        u4_sll_454_ML_int_6__92_) );
  MUX2_X2 u4_sll_454_M1_5_93 ( .A(u4_sll_454_ML_int_5__93_), .B(
        u4_sll_454_ML_int_5__61_), .S(u4_sll_454_n43), .Z(
        u4_sll_454_ML_int_6__93_) );
  MUX2_X2 u4_sll_454_M1_5_94 ( .A(u4_sll_454_ML_int_5__94_), .B(
        u4_sll_454_ML_int_5__62_), .S(u4_sll_454_n43), .Z(
        u4_sll_454_ML_int_6__94_) );
  MUX2_X2 u4_sll_454_M1_5_95 ( .A(u4_sll_454_ML_int_5__95_), .B(
        u4_sll_454_ML_int_5__63_), .S(u4_sll_454_n43), .Z(
        u4_sll_454_ML_int_6__95_) );
  MUX2_X2 u4_sll_454_M1_5_96 ( .A(u4_sll_454_ML_int_5__96_), .B(
        u4_sll_454_ML_int_5__64_), .S(u4_sll_454_n43), .Z(
        u4_sll_454_ML_int_6__96_) );
  MUX2_X2 u4_sll_454_M1_5_97 ( .A(u4_sll_454_ML_int_5__97_), .B(
        u4_sll_454_ML_int_5__65_), .S(u4_sll_454_n43), .Z(
        u4_sll_454_ML_int_6__97_) );
  MUX2_X2 u4_sll_454_M1_5_98 ( .A(u4_sll_454_ML_int_5__98_), .B(
        u4_sll_454_ML_int_5__66_), .S(u4_sll_454_n43), .Z(
        u4_sll_454_ML_int_6__98_) );
  MUX2_X2 u4_sll_454_M1_5_99 ( .A(u4_sll_454_ML_int_5__99_), .B(
        u4_sll_454_ML_int_5__67_), .S(u4_sll_454_n43), .Z(
        u4_sll_454_ML_int_6__99_) );
  MUX2_X2 u4_sll_454_M1_5_100 ( .A(u4_sll_454_ML_int_5__100_), .B(
        u4_sll_454_ML_int_5__68_), .S(u4_sll_454_n43), .Z(
        u4_sll_454_ML_int_6__100_) );
  MUX2_X2 u4_sll_454_M1_5_101 ( .A(u4_sll_454_ML_int_5__101_), .B(
        u4_sll_454_ML_int_5__69_), .S(u4_sll_454_n43), .Z(
        u4_sll_454_ML_int_6__101_) );
  MUX2_X2 u4_sll_454_M1_5_102 ( .A(u4_sll_454_ML_int_5__102_), .B(
        u4_sll_454_ML_int_5__70_), .S(u4_sll_454_n43), .Z(
        u4_sll_454_ML_int_6__102_) );
  MUX2_X2 u4_sll_454_M1_5_103 ( .A(u4_sll_454_ML_int_5__103_), .B(
        u4_sll_454_ML_int_5__71_), .S(u4_sll_454_n43), .Z(
        u4_sll_454_ML_int_6__103_) );
  MUX2_X2 u4_sll_454_M1_5_104 ( .A(u4_sll_454_ML_int_5__104_), .B(
        u4_sll_454_ML_int_5__72_), .S(u4_sll_454_n43), .Z(
        u4_sll_454_ML_int_6__104_) );
  MUX2_X2 u4_sll_454_M1_5_105 ( .A(u4_sll_454_ML_int_5__105_), .B(
        u4_sll_454_ML_int_5__73_), .S(u4_sll_454_n43), .Z(
        u4_sll_454_ML_int_6__105_) );
  MUX2_X2 u4_sll_454_M1_6_64 ( .A(u4_sll_454_ML_int_6__64_), .B(
        u4_sll_454_ML_int_6__0_), .S(u4_sll_454_n37), .Z(
        u4_sll_454_ML_int_7__64_) );
  MUX2_X2 u4_sll_454_M1_6_65 ( .A(u4_sll_454_ML_int_6__65_), .B(
        u4_sll_454_ML_int_6__1_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__65_) );
  MUX2_X2 u4_sll_454_M1_6_66 ( .A(u4_sll_454_ML_int_6__66_), .B(
        u4_sll_454_ML_int_6__2_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__66_) );
  MUX2_X2 u4_sll_454_M1_6_67 ( .A(u4_sll_454_ML_int_6__67_), .B(
        u4_sll_454_ML_int_6__3_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__67_) );
  MUX2_X2 u4_sll_454_M1_6_68 ( .A(u4_sll_454_ML_int_6__68_), .B(
        u4_sll_454_ML_int_6__4_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__68_) );
  MUX2_X2 u4_sll_454_M1_6_69 ( .A(u4_sll_454_ML_int_6__69_), .B(
        u4_sll_454_ML_int_6__5_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__69_) );
  MUX2_X2 u4_sll_454_M1_6_70 ( .A(u4_sll_454_ML_int_6__70_), .B(
        u4_sll_454_ML_int_6__6_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__70_) );
  MUX2_X2 u4_sll_454_M1_6_71 ( .A(u4_sll_454_ML_int_6__71_), .B(
        u4_sll_454_ML_int_6__7_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__71_) );
  MUX2_X2 u4_sll_454_M1_6_72 ( .A(u4_sll_454_ML_int_6__72_), .B(
        u4_sll_454_ML_int_6__8_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__72_) );
  MUX2_X2 u4_sll_454_M1_6_73 ( .A(u4_sll_454_ML_int_6__73_), .B(
        u4_sll_454_ML_int_6__9_), .S(u4_sll_454_n37), .Z(
        u4_sll_454_ML_int_7__73_) );
  MUX2_X2 u4_sll_454_M1_6_74 ( .A(u4_sll_454_ML_int_6__74_), .B(
        u4_sll_454_ML_int_6__10_), .S(u4_sll_454_n37), .Z(
        u4_sll_454_ML_int_7__74_) );
  MUX2_X2 u4_sll_454_M1_6_75 ( .A(u4_sll_454_ML_int_6__75_), .B(
        u4_sll_454_ML_int_6__11_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__75_) );
  MUX2_X2 u4_sll_454_M1_6_76 ( .A(u4_sll_454_ML_int_6__76_), .B(
        u4_sll_454_ML_int_6__12_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__76_) );
  MUX2_X2 u4_sll_454_M1_6_77 ( .A(u4_sll_454_ML_int_6__77_), .B(
        u4_sll_454_ML_int_6__13_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__77_) );
  MUX2_X2 u4_sll_454_M1_6_78 ( .A(u4_sll_454_ML_int_6__78_), .B(
        u4_sll_454_ML_int_6__14_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__78_) );
  MUX2_X2 u4_sll_454_M1_6_79 ( .A(u4_sll_454_ML_int_6__79_), .B(
        u4_sll_454_ML_int_6__15_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__79_) );
  MUX2_X2 u4_sll_454_M1_6_80 ( .A(u4_sll_454_ML_int_6__80_), .B(
        u4_sll_454_ML_int_6__16_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__80_) );
  MUX2_X2 u4_sll_454_M1_6_81 ( .A(u4_sll_454_ML_int_6__81_), .B(
        u4_sll_454_ML_int_6__17_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__81_) );
  MUX2_X2 u4_sll_454_M1_6_82 ( .A(u4_sll_454_ML_int_6__82_), .B(
        u4_sll_454_ML_int_6__18_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__82_) );
  MUX2_X2 u4_sll_454_M1_6_83 ( .A(u4_sll_454_ML_int_6__83_), .B(
        u4_sll_454_ML_int_6__19_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__83_) );
  MUX2_X2 u4_sll_454_M1_6_84 ( .A(u4_sll_454_ML_int_6__84_), .B(
        u4_sll_454_ML_int_6__20_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__84_) );
  MUX2_X2 u4_sll_454_M1_6_85 ( .A(u4_sll_454_ML_int_6__85_), .B(
        u4_sll_454_ML_int_6__21_), .S(u4_sll_454_n37), .Z(
        u4_sll_454_ML_int_7__85_) );
  MUX2_X2 u4_sll_454_M1_6_86 ( .A(u4_sll_454_ML_int_6__86_), .B(
        u4_sll_454_ML_int_6__22_), .S(u4_sll_454_n37), .Z(
        u4_sll_454_ML_int_7__86_) );
  MUX2_X2 u4_sll_454_M1_6_87 ( .A(u4_sll_454_ML_int_6__87_), .B(
        u4_sll_454_ML_int_6__23_), .S(u4_sll_454_n37), .Z(
        u4_sll_454_ML_int_7__87_) );
  MUX2_X2 u4_sll_454_M1_6_88 ( .A(u4_sll_454_ML_int_6__88_), .B(
        u4_sll_454_ML_int_6__24_), .S(u4_sll_454_n37), .Z(
        u4_sll_454_ML_int_7__88_) );
  MUX2_X2 u4_sll_454_M1_6_89 ( .A(u4_sll_454_ML_int_6__89_), .B(
        u4_sll_454_ML_int_6__25_), .S(u4_sll_454_n37), .Z(
        u4_sll_454_ML_int_7__89_) );
  MUX2_X2 u4_sll_454_M1_6_90 ( .A(u4_sll_454_ML_int_6__90_), .B(
        u4_sll_454_ML_int_6__26_), .S(u4_sll_454_n37), .Z(
        u4_sll_454_ML_int_7__90_) );
  MUX2_X2 u4_sll_454_M1_6_91 ( .A(u4_sll_454_ML_int_6__91_), .B(
        u4_sll_454_ML_int_6__27_), .S(u4_sll_454_n37), .Z(
        u4_sll_454_ML_int_7__91_) );
  MUX2_X2 u4_sll_454_M1_6_92 ( .A(u4_sll_454_ML_int_6__92_), .B(
        u4_sll_454_ML_int_6__28_), .S(u4_sll_454_n37), .Z(
        u4_sll_454_ML_int_7__92_) );
  MUX2_X2 u4_sll_454_M1_6_93 ( .A(u4_sll_454_ML_int_6__93_), .B(
        u4_sll_454_ML_int_6__29_), .S(u4_sll_454_n37), .Z(
        u4_sll_454_ML_int_7__93_) );
  MUX2_X2 u4_sll_454_M1_6_94 ( .A(u4_sll_454_ML_int_6__94_), .B(
        u4_sll_454_ML_int_6__30_), .S(u4_sll_454_n37), .Z(
        u4_sll_454_ML_int_7__94_) );
  MUX2_X2 u4_sll_454_M1_6_95 ( .A(u4_sll_454_ML_int_6__95_), .B(
        u4_sll_454_ML_int_6__31_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__95_) );
  MUX2_X2 u4_sll_454_M1_6_96 ( .A(u4_sll_454_ML_int_6__96_), .B(
        u4_sll_454_ML_int_6__32_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__96_) );
  MUX2_X2 u4_sll_454_M1_6_97 ( .A(u4_sll_454_ML_int_6__97_), .B(
        u4_sll_454_ML_int_6__33_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__97_) );
  MUX2_X2 u4_sll_454_M1_6_98 ( .A(u4_sll_454_ML_int_6__98_), .B(
        u4_sll_454_ML_int_6__34_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__98_) );
  MUX2_X2 u4_sll_454_M1_6_99 ( .A(u4_sll_454_ML_int_6__99_), .B(
        u4_sll_454_ML_int_6__35_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__99_) );
  MUX2_X2 u4_sll_454_M1_6_100 ( .A(u4_sll_454_ML_int_6__100_), .B(
        u4_sll_454_ML_int_6__36_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__100_) );
  MUX2_X2 u4_sll_454_M1_6_101 ( .A(u4_sll_454_ML_int_6__101_), .B(
        u4_sll_454_ML_int_6__37_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__101_) );
  MUX2_X2 u4_sll_454_M1_6_102 ( .A(u4_sll_454_ML_int_6__102_), .B(
        u4_sll_454_ML_int_6__38_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__102_) );
  MUX2_X2 u4_sll_454_M1_6_103 ( .A(u4_sll_454_ML_int_6__103_), .B(
        u4_sll_454_ML_int_6__39_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__103_) );
  MUX2_X2 u4_sll_454_M1_6_104 ( .A(u4_sll_454_ML_int_6__104_), .B(
        u4_sll_454_ML_int_6__40_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__104_) );
  MUX2_X2 u4_sll_454_M1_6_105 ( .A(u4_sll_454_ML_int_6__105_), .B(
        u4_sll_454_ML_int_6__41_), .S(u4_sll_454_n38), .Z(
        u4_sll_454_ML_int_7__105_) );
  NOR2_X1 u4_srl_453_U987 ( .A1(u4_shift_right[1]), .A2(u4_shift_right[7]), 
        .ZN(u4_srl_453_n878) );
  INV_X1 u4_srl_453_U986 ( .A(u4_shift_right[0]), .ZN(u4_srl_453_n879) );
  AOI22_X1 u4_srl_453_U985 ( .A1(fract_denorm[71]), .A2(u4_srl_453_n42), .B1(
        fract_denorm[70]), .B2(u4_srl_453_n47), .ZN(u4_srl_453_n877) );
  OAI221_X1 u4_srl_453_U984 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n109), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n108), .A(u4_srl_453_n877), .ZN(
        u4_srl_453_n504) );
  INV_X1 u4_srl_453_U983 ( .A(u4_srl_453_n504), .ZN(u4_srl_453_n599) );
  NOR2_X1 u4_srl_453_U982 ( .A1(u4_shift_right[3]), .A2(u4_shift_right[7]), 
        .ZN(u4_srl_453_n833) );
  INV_X1 u4_srl_453_U981 ( .A(u4_srl_453_n833), .ZN(u4_srl_453_n728) );
  INV_X1 u4_srl_453_U980 ( .A(u4_shift_right[2]), .ZN(u4_srl_453_n834) );
  NOR2_X1 u4_srl_453_U979 ( .A1(u4_srl_453_n728), .A2(u4_srl_453_n834), .ZN(
        u4_srl_453_n393) );
  AOI22_X1 u4_srl_453_U978 ( .A1(fract_denorm[67]), .A2(u4_srl_453_n42), .B1(
        fract_denorm[66]), .B2(u4_srl_453_n47), .ZN(u4_srl_453_n876) );
  OAI221_X1 u4_srl_453_U977 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n105), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n104), .A(u4_srl_453_n876), .ZN(
        u4_srl_453_n505) );
  INV_X1 u4_srl_453_U976 ( .A(u4_srl_453_n505), .ZN(u4_srl_453_n746) );
  NOR2_X1 u4_srl_453_U975 ( .A1(u4_srl_453_n728), .A2(u4_shift_right[2]), .ZN(
        u4_srl_453_n409) );
  NOR2_X1 u4_srl_453_U974 ( .A1(u4_srl_453_n834), .A2(u4_srl_453_n833), .ZN(
        u4_srl_453_n394) );
  AOI22_X1 u4_srl_453_U973 ( .A1(fract_denorm[79]), .A2(u4_srl_453_n43), .B1(
        fract_denorm[78]), .B2(u4_srl_453_n49), .ZN(u4_srl_453_n875) );
  OAI221_X1 u4_srl_453_U972 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n95), .C1(
        u4_srl_453_n39), .C2(u4_srl_453_n94), .A(u4_srl_453_n875), .ZN(
        u4_srl_453_n601) );
  AOI22_X1 u4_srl_453_U971 ( .A1(fract_denorm[75]), .A2(u4_srl_453_n42), .B1(
        fract_denorm[74]), .B2(u4_srl_453_n52), .ZN(u4_srl_453_n874) );
  OAI221_X1 u4_srl_453_U970 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n112), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n111), .A(u4_srl_453_n874), .ZN(
        u4_srl_453_n602) );
  AOI22_X1 u4_srl_453_U969 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n601), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n602), .ZN(u4_srl_453_n873) );
  OAI221_X1 u4_srl_453_U968 ( .B1(u4_srl_453_n599), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n746), .C2(u4_srl_453_n59), .A(u4_srl_453_n873), .ZN(
        u4_srl_453_n423) );
  NOR2_X1 u4_srl_453_U967 ( .A1(u4_shift_right[5]), .A2(u4_shift_right[7]), 
        .ZN(u4_srl_453_n266) );
  INV_X1 u4_srl_453_U966 ( .A(u4_srl_453_n238), .ZN(u4_srl_453_n400) );
  AOI22_X1 u4_srl_453_U965 ( .A1(fract_denorm[103]), .A2(u4_srl_453_n46), .B1(
        fract_denorm[102]), .B2(u4_srl_453_n52), .ZN(u4_srl_453_n872) );
  OAI221_X1 u4_srl_453_U964 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n76), .C1(
        u4_srl_453_n37), .C2(u4_srl_453_n78), .A(u4_srl_453_n872), .ZN(
        u4_srl_453_n499) );
  AOI22_X1 u4_srl_453_U963 ( .A1(u4_srl_453_n41), .A2(fract_denorm[104]), .B1(
        u4_srl_453_n35), .B2(n4652), .ZN(u4_srl_453_n244) );
  INV_X1 u4_srl_453_U962 ( .A(u4_srl_453_n244), .ZN(u4_srl_453_n380) );
  AOI22_X1 u4_srl_453_U961 ( .A1(fract_denorm[99]), .A2(u4_srl_453_n46), .B1(
        fract_denorm[98]), .B2(u4_srl_453_n52), .ZN(u4_srl_453_n871) );
  OAI221_X1 u4_srl_453_U960 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n72), .C1(
        u4_srl_453_n40), .C2(u4_srl_453_n71), .A(u4_srl_453_n871), .ZN(
        u4_srl_453_n500) );
  AOI222_X1 u4_srl_453_U959 ( .A1(u4_srl_453_n499), .A2(u4_srl_453_n15), .B1(
        u4_srl_453_n380), .B2(u4_srl_453_n25), .C1(u4_srl_453_n500), .C2(
        u4_srl_453_n56), .ZN(u4_srl_453_n184) );
  INV_X1 u4_srl_453_U958 ( .A(u4_srl_453_n184), .ZN(u4_srl_453_n346) );
  NOR2_X1 u4_srl_453_U957 ( .A1(u4_shift_right[4]), .A2(u4_srl_453_n266), .ZN(
        u4_srl_453_n336) );
  AOI22_X1 u4_srl_453_U956 ( .A1(fract_denorm[87]), .A2(u4_srl_453_n42), .B1(
        fract_denorm[86]), .B2(u4_srl_453_n52), .ZN(u4_srl_453_n870) );
  OAI221_X1 u4_srl_453_U955 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n88), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n87), .A(u4_srl_453_n870), .ZN(
        u4_srl_453_n494) );
  INV_X1 u4_srl_453_U954 ( .A(u4_srl_453_n494), .ZN(u4_srl_453_n603) );
  AOI22_X1 u4_srl_453_U953 ( .A1(fract_denorm[83]), .A2(u4_srl_453_n42), .B1(
        fract_denorm[82]), .B2(u4_srl_453_n52), .ZN(u4_srl_453_n869) );
  OAI221_X1 u4_srl_453_U952 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n98), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n97), .A(u4_srl_453_n869), .ZN(
        u4_srl_453_n495) );
  INV_X1 u4_srl_453_U951 ( .A(u4_srl_453_n495), .ZN(u4_srl_453_n748) );
  AOI22_X1 u4_srl_453_U950 ( .A1(fract_denorm[95]), .A2(u4_srl_453_n46), .B1(
        fract_denorm[94]), .B2(u4_srl_453_n52), .ZN(u4_srl_453_n868) );
  OAI221_X1 u4_srl_453_U949 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n69), .C1(
        u4_srl_453_n39), .C2(u4_srl_453_n68), .A(u4_srl_453_n868), .ZN(
        u4_srl_453_n605) );
  AOI22_X1 u4_srl_453_U948 ( .A1(fract_denorm[91]), .A2(u4_srl_453_n46), .B1(
        fract_denorm[90]), .B2(u4_srl_453_n52), .ZN(u4_srl_453_n867) );
  OAI221_X1 u4_srl_453_U947 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n91), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n90), .A(u4_srl_453_n867), .ZN(
        u4_srl_453_n606) );
  AOI22_X1 u4_srl_453_U946 ( .A1(u4_srl_453_n23), .A2(u4_srl_453_n605), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n606), .ZN(u4_srl_453_n866) );
  OAI221_X1 u4_srl_453_U945 ( .B1(u4_srl_453_n603), .B2(u4_srl_453_n19), .C1(
        u4_srl_453_n748), .C2(u4_srl_453_n58), .A(u4_srl_453_n866), .ZN(
        u4_srl_453_n347) );
  INV_X1 u4_srl_453_U944 ( .A(u4_srl_453_n242), .ZN(u4_srl_453_n401) );
  AOI222_X1 u4_srl_453_U943 ( .A1(u4_srl_453_n423), .A2(u4_srl_453_n400), .B1(
        u4_srl_453_n346), .B2(u4_srl_453_n336), .C1(u4_srl_453_n347), .C2(
        u4_srl_453_n401), .ZN(u4_srl_453_n272) );
  NOR2_X1 u4_srl_453_U942 ( .A1(u4_shift_right[6]), .A2(u4_shift_right[7]), 
        .ZN(u4_srl_453_n859) );
  NOR2_X1 u4_srl_453_U941 ( .A1(u4_srl_453_n859), .A2(u4_shift_right[8]), .ZN(
        u4_srl_453_n376) );
  AOI22_X1 u4_srl_453_U940 ( .A1(fract_denorm[55]), .A2(u4_srl_453_n42), .B1(
        fract_denorm[54]), .B2(u4_srl_453_n52), .ZN(u4_srl_453_n865) );
  OAI221_X1 u4_srl_453_U939 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n81), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n114), .A(u4_srl_453_n865), .ZN(
        u4_srl_453_n517) );
  AOI22_X1 u4_srl_453_U938 ( .A1(fract_denorm[51]), .A2(u4_srl_453_n43), .B1(
        fract_denorm[50]), .B2(u4_srl_453_n52), .ZN(u4_srl_453_n864) );
  OAI221_X1 u4_srl_453_U937 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n80), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n125), .A(u4_srl_453_n864), .ZN(
        u4_srl_453_n518) );
  AOI22_X1 u4_srl_453_U936 ( .A1(fract_denorm[63]), .A2(u4_srl_453_n42), .B1(
        fract_denorm[62]), .B2(u4_srl_453_n52), .ZN(u4_srl_453_n863) );
  OAI221_X1 u4_srl_453_U935 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n102), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n101), .A(u4_srl_453_n863), .ZN(
        u4_srl_453_n609) );
  AOI22_X1 u4_srl_453_U934 ( .A1(fract_denorm[59]), .A2(u4_srl_453_n43), .B1(
        fract_denorm[58]), .B2(u4_srl_453_n52), .ZN(u4_srl_453_n862) );
  OAI221_X1 u4_srl_453_U933 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n84), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n83), .A(u4_srl_453_n862), .ZN(
        u4_srl_453_n506) );
  AOI22_X1 u4_srl_453_U932 ( .A1(u4_srl_453_n23), .A2(u4_srl_453_n609), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n506), .ZN(u4_srl_453_n861) );
  INV_X1 u4_srl_453_U931 ( .A(u4_srl_453_n861), .ZN(u4_srl_453_n860) );
  AOI221_X1 u4_srl_453_U930 ( .B1(u4_srl_453_n517), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n518), .C2(u4_srl_453_n56), .A(u4_srl_453_n860), .ZN(
        u4_srl_453_n344) );
  NOR2_X1 u4_srl_453_U929 ( .A1(u4_srl_453_n174), .A2(u4_srl_453_n266), .ZN(
        u4_srl_453_n801) );
  INV_X1 u4_srl_453_U928 ( .A(u4_shift_right[8]), .ZN(u4_srl_453_n858) );
  NAND2_X1 u4_srl_453_U927 ( .A1(u4_srl_453_n801), .A2(u4_srl_453_n858), .ZN(
        u4_srl_453_n299) );
  NOR2_X1 u4_srl_453_U926 ( .A1(u4_srl_453_n299), .A2(u4_srl_453_n392), .ZN(
        u4_srl_453_n312) );
  AOI22_X1 u4_srl_453_U925 ( .A1(n6439), .A2(u4_srl_453_n45), .B1(n6436), .B2(
        u4_srl_453_n52), .ZN(u4_srl_453_n857) );
  OAI221_X1 u4_srl_453_U924 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n149), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n148), .A(u4_srl_453_n857), .ZN(
        u4_srl_453_n510) );
  AOI22_X1 u4_srl_453_U923 ( .A1(n6433), .A2(u4_srl_453_n45), .B1(n6440), .B2(
        u4_srl_453_n51), .ZN(u4_srl_453_n856) );
  OAI221_X1 u4_srl_453_U922 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n145), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n144), .A(u4_srl_453_n856), .ZN(
        u4_srl_453_n511) );
  AOI22_X1 u4_srl_453_U921 ( .A1(n6410), .A2(u4_srl_453_n45), .B1(n6408), .B2(
        u4_srl_453_n51), .ZN(u4_srl_453_n855) );
  OAI221_X1 u4_srl_453_U920 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n123), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n122), .A(u4_srl_453_n855), .ZN(
        u4_srl_453_n513) );
  AOI22_X1 u4_srl_453_U919 ( .A1(n6405), .A2(u4_srl_453_n45), .B1(n6445), .B2(
        u4_srl_453_n51), .ZN(u4_srl_453_n854) );
  OAI221_X1 u4_srl_453_U918 ( .B1(u4_srl_453_n32), .B2(u4_srl_453_n152), .C1(
        u4_srl_453_n40), .C2(u4_srl_453_n151), .A(u4_srl_453_n854), .ZN(
        u4_srl_453_n514) );
  AOI22_X1 u4_srl_453_U917 ( .A1(u4_srl_453_n23), .A2(u4_srl_453_n513), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n514), .ZN(u4_srl_453_n853) );
  INV_X1 u4_srl_453_U916 ( .A(u4_srl_453_n853), .ZN(u4_srl_453_n852) );
  AOI221_X1 u4_srl_453_U915 ( .B1(u4_srl_453_n510), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n511), .C2(u4_srl_453_n409), .A(u4_srl_453_n852), .ZN(
        u4_srl_453_n421) );
  INV_X1 u4_srl_453_U914 ( .A(u4_srl_453_n421), .ZN(u4_srl_453_n837) );
  NAND2_X1 u4_srl_453_U913 ( .A1(u4_srl_453_n210), .A2(u4_srl_453_n266), .ZN(
        u4_srl_453_n204) );
  INV_X1 u4_srl_453_U912 ( .A(u4_srl_453_n204), .ZN(u4_srl_453_n386) );
  OAI22_X1 u4_srl_453_U911 ( .A1(u4_srl_453_n54), .A2(u4_srl_453_n60), .B1(
        u4_srl_453_n1), .B2(u4_srl_453_n61), .ZN(u4_srl_453_n851) );
  AOI221_X1 u4_srl_453_U910 ( .B1(n6344), .B2(u4_srl_453_n35), .C1(n6446), 
        .C2(u4_srl_453_n41), .A(u4_srl_453_n851), .ZN(u4_srl_453_n839) );
  NAND2_X1 u4_srl_453_U909 ( .A1(u4_srl_453_n409), .A2(u4_srl_453_n392), .ZN(
        u4_srl_453_n265) );
  OAI22_X1 u4_srl_453_U908 ( .A1(u4_srl_453_n139), .A2(u4_srl_453_n1), .B1(
        u4_srl_453_n136), .B2(u4_srl_453_n54), .ZN(u4_srl_453_n850) );
  AOI221_X1 u4_srl_453_U907 ( .B1(u4_srl_453_n35), .B2(n6421), .C1(
        u4_srl_453_n41), .C2(n6420), .A(u4_srl_453_n850), .ZN(u4_srl_453_n197)
         );
  AOI22_X1 u4_srl_453_U906 ( .A1(n6419), .A2(u4_srl_453_n45), .B1(n6442), .B2(
        u4_srl_453_n51), .ZN(u4_srl_453_n849) );
  OAI221_X1 u4_srl_453_U905 ( .B1(u4_srl_453_n32), .B2(u4_srl_453_n132), .C1(
        u4_srl_453_n40), .C2(u4_srl_453_n131), .A(u4_srl_453_n849), .ZN(
        u4_srl_453_n327) );
  INV_X1 u4_srl_453_U904 ( .A(u4_srl_453_n327), .ZN(u4_srl_453_n196) );
  AOI22_X1 u4_srl_453_U903 ( .A1(n6432), .A2(u4_srl_453_n45), .B1(n6429), .B2(
        u4_srl_453_n51), .ZN(u4_srl_453_n848) );
  OAI221_X1 u4_srl_453_U902 ( .B1(u4_srl_453_n32), .B2(u4_srl_453_n142), .C1(
        u4_srl_453_n40), .C2(u4_srl_453_n141), .A(u4_srl_453_n848), .ZN(
        u4_srl_453_n512) );
  AOI22_X1 u4_srl_453_U901 ( .A1(n6426), .A2(u4_srl_453_n45), .B1(n6441), .B2(
        u4_srl_453_n51), .ZN(u4_srl_453_n847) );
  OAI221_X1 u4_srl_453_U900 ( .B1(u4_srl_453_n32), .B2(u4_srl_453_n138), .C1(
        u4_srl_453_n137), .C2(u4_srl_453_n36), .A(u4_srl_453_n847), .ZN(
        u4_srl_453_n741) );
  AOI22_X1 u4_srl_453_U899 ( .A1(u4_srl_453_n23), .A2(u4_srl_453_n512), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n741), .ZN(u4_srl_453_n846) );
  OAI221_X1 u4_srl_453_U898 ( .B1(u4_srl_453_n197), .B2(u4_srl_453_n19), .C1(
        u4_srl_453_n196), .C2(u4_srl_453_n58), .A(u4_srl_453_n846), .ZN(
        u4_srl_453_n845) );
  INV_X1 u4_srl_453_U897 ( .A(u4_srl_453_n845), .ZN(u4_srl_453_n673) );
  AOI22_X1 u4_srl_453_U896 ( .A1(n6350), .A2(u4_srl_453_n45), .B1(n6349), .B2(
        u4_srl_453_n51), .ZN(u4_srl_453_n844) );
  OAI221_X1 u4_srl_453_U895 ( .B1(u4_srl_453_n32), .B2(u4_srl_453_n63), .C1(
        u4_srl_453_n40), .C2(u4_srl_453_n62), .A(u4_srl_453_n844), .ZN(
        u4_srl_453_n330) );
  AOI22_X1 u4_srl_453_U894 ( .A1(n6418), .A2(u4_srl_453_n45), .B1(n6415), .B2(
        u4_srl_453_n51), .ZN(u4_srl_453_n843) );
  OAI221_X1 u4_srl_453_U893 ( .B1(u4_srl_453_n32), .B2(u4_srl_453_n129), .C1(
        u4_srl_453_n40), .C2(u4_srl_453_n128), .A(u4_srl_453_n843), .ZN(
        u4_srl_453_n193) );
  AOI22_X1 u4_srl_453_U892 ( .A1(n6411), .A2(u4_srl_453_n45), .B1(n6443), .B2(
        u4_srl_453_n51), .ZN(u4_srl_453_n842) );
  OAI221_X1 u4_srl_453_U891 ( .B1(u4_srl_453_n32), .B2(u4_srl_453_n158), .C1(
        u4_srl_453_n40), .C2(u4_srl_453_n66), .A(u4_srl_453_n842), .ZN(
        u4_srl_453_n194) );
  AOI222_X1 u4_srl_453_U890 ( .A1(u4_srl_453_n15), .A2(u4_srl_453_n330), .B1(
        u4_srl_453_n21), .B2(u4_srl_453_n193), .C1(u4_srl_453_n25), .C2(
        u4_srl_453_n194), .ZN(u4_srl_453_n841) );
  MUX2_X1 u4_srl_453_U889 ( .A(u4_srl_453_n673), .B(u4_srl_453_n841), .S(
        u4_srl_453_n392), .Z(u4_srl_453_n840) );
  OAI21_X1 u4_srl_453_U888 ( .B1(u4_srl_453_n839), .B2(u4_srl_453_n265), .A(
        u4_srl_453_n840), .ZN(u4_srl_453_n838) );
  AOI22_X1 u4_srl_453_U887 ( .A1(u4_srl_453_n14), .A2(u4_srl_453_n837), .B1(
        u4_srl_453_n386), .B2(u4_srl_453_n838), .ZN(u4_srl_453_n836) );
  OAI221_X1 u4_srl_453_U886 ( .B1(u4_srl_453_n272), .B2(u4_srl_453_n383), .C1(
        u4_srl_453_n344), .C2(u4_srl_453_n11), .A(u4_srl_453_n836), .ZN(
        u4_N5906) );
  AOI22_X1 u4_srl_453_U885 ( .A1(u4_srl_453_n499), .A2(u4_srl_453_n409), .B1(
        u4_srl_453_n380), .B2(u4_srl_453_n16), .ZN(u4_srl_453_n334) );
  NAND2_X1 u4_srl_453_U884 ( .A1(u4_srl_453_n386), .A2(u4_srl_453_n392), .ZN(
        u4_srl_453_n181) );
  NOR2_X1 u4_srl_453_U883 ( .A1(u4_srl_453_n334), .A2(u4_srl_453_n8), .ZN(
        u4_N6006) );
  NAND2_X1 u4_srl_453_U882 ( .A1(n4652), .A2(u4_srl_453_n41), .ZN(
        u4_srl_453_n240) );
  INV_X1 u4_srl_453_U881 ( .A(u4_srl_453_n240), .ZN(u4_srl_453_n665) );
  AOI22_X1 u4_srl_453_U880 ( .A1(fract_denorm[104]), .A2(u4_srl_453_n45), .B1(
        fract_denorm[103]), .B2(u4_srl_453_n51), .ZN(u4_srl_453_n835) );
  OAI221_X1 u4_srl_453_U879 ( .B1(u4_srl_453_n32), .B2(u4_srl_453_n77), .C1(
        u4_srl_453_n40), .C2(u4_srl_453_n76), .A(u4_srl_453_n835), .ZN(
        u4_srl_453_n469) );
  MUX2_X1 u4_srl_453_U878 ( .A(u4_srl_453_n665), .B(u4_srl_453_n469), .S(
        u4_srl_453_n834), .Z(u4_srl_453_n729) );
  NAND2_X1 u4_srl_453_U877 ( .A1(u4_srl_453_n833), .A2(u4_srl_453_n729), .ZN(
        u4_srl_453_n292) );
  NOR2_X1 u4_srl_453_U876 ( .A1(u4_srl_453_n181), .A2(u4_srl_453_n292), .ZN(
        u4_N6007) );
  AOI22_X1 u4_srl_453_U875 ( .A1(n4652), .A2(u4_srl_453_n45), .B1(
        fract_denorm[104]), .B2(u4_srl_453_n51), .ZN(u4_srl_453_n832) );
  INV_X1 u4_srl_453_U874 ( .A(u4_srl_453_n832), .ZN(u4_srl_453_n831) );
  AOI221_X1 u4_srl_453_U873 ( .B1(u4_srl_453_n35), .B2(fract_denorm[103]), 
        .C1(u4_srl_453_n41), .C2(fract_denorm[102]), .A(u4_srl_453_n831), .ZN(
        u4_srl_453_n263) );
  OR2_X1 u4_srl_453_U872 ( .A1(u4_srl_453_n181), .A2(u4_srl_453_n59), .ZN(
        u4_srl_453_n830) );
  NOR2_X1 u4_srl_453_U871 ( .A1(u4_srl_453_n263), .A2(u4_srl_453_n830), .ZN(
        u4_N6008) );
  AOI222_X1 u4_srl_453_U870 ( .A1(u4_srl_453_n35), .A2(fract_denorm[104]), 
        .B1(u4_srl_453_n47), .B2(n4652), .C1(u4_srl_453_n41), .C2(
        fract_denorm[103]), .ZN(u4_srl_453_n247) );
  NOR2_X1 u4_srl_453_U869 ( .A1(u4_srl_453_n247), .A2(u4_srl_453_n830), .ZN(
        u4_N6009) );
  NOR2_X1 u4_srl_453_U868 ( .A1(u4_srl_453_n244), .A2(u4_srl_453_n830), .ZN(
        u4_N6010) );
  NOR3_X1 u4_srl_453_U867 ( .A1(u4_srl_453_n58), .A2(u4_srl_453_n238), .A3(
        u4_srl_453_n240), .ZN(u4_srl_453_n375) );
  AND2_X1 u4_srl_453_U866 ( .A1(u4_srl_453_n210), .A2(u4_srl_453_n375), .ZN(
        u4_N6011) );
  AOI22_X1 u4_srl_453_U865 ( .A1(n6431), .A2(u4_srl_453_n43), .B1(n6430), .B2(
        u4_srl_453_n51), .ZN(u4_srl_453_n829) );
  OAI221_X1 u4_srl_453_U864 ( .B1(u4_srl_453_n32), .B2(u4_srl_453_n146), .C1(
        u4_srl_453_n40), .C2(u4_srl_453_n143), .A(u4_srl_453_n829), .ZN(
        u4_srl_453_n574) );
  AOI22_X1 u4_srl_453_U863 ( .A1(n6428), .A2(u4_srl_453_n42), .B1(n6427), .B2(
        u4_srl_453_n50), .ZN(u4_srl_453_n828) );
  OAI221_X1 u4_srl_453_U862 ( .B1(u4_srl_453_n32), .B2(u4_srl_453_n140), .C1(
        u4_srl_453_n40), .C2(u4_srl_453_n155), .A(u4_srl_453_n828), .ZN(
        u4_srl_453_n655) );
  AOI22_X1 u4_srl_453_U861 ( .A1(n6438), .A2(u4_srl_453_n43), .B1(n6437), .B2(
        u4_srl_453_n50), .ZN(u4_srl_453_n827) );
  OAI221_X1 u4_srl_453_U860 ( .B1(u4_srl_453_n32), .B2(u4_srl_453_n153), .C1(
        u4_srl_453_n40), .C2(u4_srl_453_n150), .A(u4_srl_453_n827), .ZN(
        u4_srl_453_n576) );
  AOI22_X1 u4_srl_453_U859 ( .A1(n6435), .A2(u4_srl_453_n42), .B1(n6434), .B2(
        u4_srl_453_n50), .ZN(u4_srl_453_n826) );
  OAI221_X1 u4_srl_453_U858 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n147), .C1(
        u4_srl_453_n40), .C2(u4_srl_453_n154), .A(u4_srl_453_n826), .ZN(
        u4_srl_453_n573) );
  AOI22_X1 u4_srl_453_U857 ( .A1(u4_srl_453_n23), .A2(u4_srl_453_n576), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n573), .ZN(u4_srl_453_n825) );
  INV_X1 u4_srl_453_U856 ( .A(u4_srl_453_n825), .ZN(u4_srl_453_n824) );
  AOI221_X1 u4_srl_453_U855 ( .B1(u4_srl_453_n574), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n655), .C2(u4_srl_453_n409), .A(u4_srl_453_n824), .ZN(
        u4_srl_453_n452) );
  INV_X1 u4_srl_453_U854 ( .A(u4_srl_453_n452), .ZN(u4_srl_453_n799) );
  AOI22_X1 u4_srl_453_U853 ( .A1(fract_denorm[97]), .A2(u4_srl_453_n46), .B1(
        fract_denorm[96]), .B2(u4_srl_453_n50), .ZN(u4_srl_453_n823) );
  OAI221_X1 u4_srl_453_U852 ( .B1(u4_srl_453_n2), .B2(u4_srl_453_n73), .C1(
        u4_srl_453_n6), .C2(u4_srl_453_n70), .A(u4_srl_453_n823), .ZN(
        u4_srl_453_n563) );
  AOI22_X1 u4_srl_453_U851 ( .A1(fract_denorm[93]), .A2(u4_srl_453_n44), .B1(
        fract_denorm[92]), .B2(u4_srl_453_n50), .ZN(u4_srl_453_n822) );
  OAI221_X1 u4_srl_453_U850 ( .B1(u4_srl_453_n32), .B2(u4_srl_453_n67), .C1(
        u4_srl_453_n40), .C2(u4_srl_453_n74), .A(u4_srl_453_n822), .ZN(
        u4_srl_453_n558) );
  INV_X1 u4_srl_453_U849 ( .A(u4_srl_453_n263), .ZN(u4_srl_453_n406) );
  AOI22_X1 u4_srl_453_U848 ( .A1(fract_denorm[101]), .A2(u4_srl_453_n46), .B1(
        fract_denorm[100]), .B2(u4_srl_453_n50), .ZN(u4_srl_453_n821) );
  OAI221_X1 u4_srl_453_U847 ( .B1(u4_srl_453_n2), .B2(u4_srl_453_n75), .C1(
        u4_srl_453_n6), .C2(u4_srl_453_n79), .A(u4_srl_453_n821), .ZN(
        u4_srl_453_n562) );
  AOI22_X1 u4_srl_453_U846 ( .A1(u4_srl_453_n23), .A2(u4_srl_453_n406), .B1(
        u4_srl_453_n28), .B2(u4_srl_453_n562), .ZN(u4_srl_453_n820) );
  INV_X1 u4_srl_453_U845 ( .A(u4_srl_453_n820), .ZN(u4_srl_453_n819) );
  AOI221_X1 u4_srl_453_U844 ( .B1(u4_srl_453_n563), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n558), .C2(u4_srl_453_n57), .A(u4_srl_453_n819), .ZN(
        u4_srl_453_n190) );
  AOI22_X1 u4_srl_453_U843 ( .A1(fract_denorm[81]), .A2(u4_srl_453_n43), .B1(
        fract_denorm[80]), .B2(u4_srl_453_n50), .ZN(u4_srl_453_n818) );
  OAI221_X1 u4_srl_453_U842 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n99), .C1(
        u4_srl_453_n37), .C2(u4_srl_453_n96), .A(u4_srl_453_n818), .ZN(
        u4_srl_453_n557) );
  INV_X1 u4_srl_453_U841 ( .A(u4_srl_453_n557), .ZN(u4_srl_453_n698) );
  AOI22_X1 u4_srl_453_U840 ( .A1(fract_denorm[77]), .A2(u4_srl_453_n45), .B1(
        fract_denorm[76]), .B2(u4_srl_453_n50), .ZN(u4_srl_453_n817) );
  OAI221_X1 u4_srl_453_U839 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n93), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n118), .A(u4_srl_453_n817), .ZN(
        u4_srl_453_n645) );
  INV_X1 u4_srl_453_U838 ( .A(u4_srl_453_n645), .ZN(u4_srl_453_n553) );
  AOI22_X1 u4_srl_453_U837 ( .A1(fract_denorm[89]), .A2(u4_srl_453_n46), .B1(
        fract_denorm[88]), .B2(u4_srl_453_n50), .ZN(u4_srl_453_n816) );
  OAI221_X1 u4_srl_453_U836 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n92), .C1(
        u4_srl_453_n39), .C2(u4_srl_453_n89), .A(u4_srl_453_n816), .ZN(
        u4_srl_453_n559) );
  AOI22_X1 u4_srl_453_U835 ( .A1(fract_denorm[85]), .A2(u4_srl_453_n42), .B1(
        fract_denorm[84]), .B2(u4_srl_453_n50), .ZN(u4_srl_453_n815) );
  OAI221_X1 u4_srl_453_U834 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n86), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n117), .A(u4_srl_453_n815), .ZN(
        u4_srl_453_n556) );
  AOI22_X1 u4_srl_453_U833 ( .A1(u4_srl_453_n23), .A2(u4_srl_453_n559), .B1(
        u4_srl_453_n28), .B2(u4_srl_453_n556), .ZN(u4_srl_453_n814) );
  OAI221_X1 u4_srl_453_U832 ( .B1(u4_srl_453_n698), .B2(u4_srl_453_n19), .C1(
        u4_srl_453_n553), .C2(u4_srl_453_n59), .A(u4_srl_453_n814), .ZN(
        u4_srl_453_n371) );
  INV_X1 u4_srl_453_U831 ( .A(u4_srl_453_n371), .ZN(u4_srl_453_n297) );
  OAI22_X1 u4_srl_453_U830 ( .A1(u4_srl_453_n190), .A2(u4_srl_453_n242), .B1(
        u4_srl_453_n297), .B2(u4_srl_453_n238), .ZN(u4_srl_453_n236) );
  AOI22_X1 u4_srl_453_U829 ( .A1(fract_denorm[65]), .A2(u4_srl_453_n43), .B1(
        fract_denorm[64]), .B2(u4_srl_453_n50), .ZN(u4_srl_453_n813) );
  OAI221_X1 u4_srl_453_U828 ( .B1(u4_srl_453_n32), .B2(u4_srl_453_n106), .C1(
        u4_srl_453_n40), .C2(u4_srl_453_n103), .A(u4_srl_453_n813), .ZN(
        u4_srl_453_n569) );
  AOI22_X1 u4_srl_453_U827 ( .A1(fract_denorm[61]), .A2(u4_srl_453_n44), .B1(
        fract_denorm[60]), .B2(u4_srl_453_n50), .ZN(u4_srl_453_n812) );
  OAI221_X1 u4_srl_453_U826 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n100), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n115), .A(u4_srl_453_n812), .ZN(
        u4_srl_453_n564) );
  AOI22_X1 u4_srl_453_U825 ( .A1(fract_denorm[73]), .A2(u4_srl_453_n44), .B1(
        fract_denorm[72]), .B2(u4_srl_453_n51), .ZN(u4_srl_453_n811) );
  OAI221_X1 u4_srl_453_U824 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n113), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n110), .A(u4_srl_453_n811), .ZN(
        u4_srl_453_n646) );
  AOI22_X1 u4_srl_453_U823 ( .A1(fract_denorm[69]), .A2(u4_srl_453_n44), .B1(
        fract_denorm[68]), .B2(u4_srl_453_n49), .ZN(u4_srl_453_n810) );
  OAI221_X1 u4_srl_453_U822 ( .B1(u4_srl_453_n31), .B2(u4_srl_453_n107), .C1(
        u4_srl_453_n39), .C2(u4_srl_453_n116), .A(u4_srl_453_n810), .ZN(
        u4_srl_453_n568) );
  AOI22_X1 u4_srl_453_U821 ( .A1(u4_srl_453_n23), .A2(u4_srl_453_n646), .B1(
        u4_srl_453_n27), .B2(u4_srl_453_n568), .ZN(u4_srl_453_n809) );
  INV_X1 u4_srl_453_U820 ( .A(u4_srl_453_n809), .ZN(u4_srl_453_n808) );
  AOI221_X1 u4_srl_453_U819 ( .B1(u4_srl_453_n569), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n564), .C2(u4_srl_453_n57), .A(u4_srl_453_n808), .ZN(
        u4_srl_453_n298) );
  AOI22_X1 u4_srl_453_U818 ( .A1(n6367), .A2(u4_srl_453_n44), .B1(n6409), .B2(
        u4_srl_453_n47), .ZN(u4_srl_453_n807) );
  OAI221_X1 u4_srl_453_U817 ( .B1(u4_srl_453_n31), .B2(u4_srl_453_n126), .C1(
        u4_srl_453_n39), .C2(u4_srl_453_n124), .A(u4_srl_453_n807), .ZN(
        u4_srl_453_n580) );
  AOI22_X1 u4_srl_453_U816 ( .A1(n6407), .A2(u4_srl_453_n44), .B1(n6406), .B2(
        u4_srl_453_n47), .ZN(u4_srl_453_n806) );
  OAI221_X1 u4_srl_453_U815 ( .B1(u4_srl_453_n31), .B2(u4_srl_453_n121), .C1(
        u4_srl_453_n39), .C2(u4_srl_453_n159), .A(u4_srl_453_n806), .ZN(
        u4_srl_453_n575) );
  AOI22_X1 u4_srl_453_U814 ( .A1(fract_denorm[57]), .A2(u4_srl_453_n44), .B1(
        fract_denorm[56]), .B2(u4_srl_453_n47), .ZN(u4_srl_453_n805) );
  OAI221_X1 u4_srl_453_U813 ( .B1(u4_srl_453_n31), .B2(u4_srl_453_n85), .C1(
        u4_srl_453_n39), .C2(u4_srl_453_n82), .A(u4_srl_453_n805), .ZN(
        u4_srl_453_n565) );
  AOI22_X1 u4_srl_453_U812 ( .A1(fract_denorm[53]), .A2(u4_srl_453_n44), .B1(
        fract_denorm[52]), .B2(u4_srl_453_n47), .ZN(u4_srl_453_n804) );
  OAI221_X1 u4_srl_453_U811 ( .B1(u4_srl_453_n31), .B2(u4_srl_453_n119), .C1(
        u4_srl_453_n39), .C2(u4_srl_453_n120), .A(u4_srl_453_n804), .ZN(
        u4_srl_453_n579) );
  AOI22_X1 u4_srl_453_U810 ( .A1(u4_srl_453_n23), .A2(u4_srl_453_n565), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n579), .ZN(u4_srl_453_n803) );
  INV_X1 u4_srl_453_U809 ( .A(u4_srl_453_n803), .ZN(u4_srl_453_n802) );
  AOI221_X1 u4_srl_453_U808 ( .B1(u4_srl_453_n580), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n575), .C2(u4_srl_453_n57), .A(u4_srl_453_n802), .ZN(
        u4_srl_453_n373) );
  OAI22_X1 u4_srl_453_U807 ( .A1(u4_srl_453_n298), .A2(u4_srl_453_n177), .B1(
        u4_srl_453_n373), .B2(u4_srl_453_n179), .ZN(u4_srl_453_n800) );
  AOI221_X1 u4_srl_453_U806 ( .B1(u4_srl_453_n171), .B2(u4_srl_453_n799), .C1(
        u4_srl_453_n236), .C2(u4_srl_453_n174), .A(u4_srl_453_n800), .ZN(
        u4_srl_453_n791) );
  NOR2_X1 u4_srl_453_U805 ( .A1(u4_srl_453_n238), .A2(u4_srl_453_n174), .ZN(
        u4_srl_453_n794) );
  AOI22_X1 u4_srl_453_U804 ( .A1(n6417), .A2(u4_srl_453_n44), .B1(n6416), .B2(
        u4_srl_453_n47), .ZN(u4_srl_453_n798) );
  OAI221_X1 u4_srl_453_U803 ( .B1(u4_srl_453_n31), .B2(u4_srl_453_n133), .C1(
        u4_srl_453_n39), .C2(u4_srl_453_n130), .A(u4_srl_453_n798), .ZN(
        u4_srl_453_n253) );
  AOI22_X1 u4_srl_453_U802 ( .A1(n6414), .A2(u4_srl_453_n44), .B1(n6413), .B2(
        u4_srl_453_n47), .ZN(u4_srl_453_n797) );
  OAI221_X1 u4_srl_453_U801 ( .B1(u4_srl_453_n31), .B2(u4_srl_453_n127), .C1(
        u4_srl_453_n39), .C2(u4_srl_453_n157), .A(u4_srl_453_n797), .ZN(
        u4_srl_453_n257) );
  AOI22_X1 u4_srl_453_U800 ( .A1(n6421), .A2(u4_srl_453_n44), .B1(n6420), .B2(
        u4_srl_453_n47), .ZN(u4_srl_453_n796) );
  OAI221_X1 u4_srl_453_U799 ( .B1(u4_srl_453_n31), .B2(u4_srl_453_n134), .C1(
        u4_srl_453_n39), .C2(u4_srl_453_n156), .A(u4_srl_453_n796), .ZN(
        u4_srl_453_n252) );
  INV_X1 u4_srl_453_U798 ( .A(u4_srl_453_n252), .ZN(u4_srl_453_n653) );
  OAI22_X1 u4_srl_453_U797 ( .A1(u4_srl_453_n138), .A2(u4_srl_453_n1), .B1(
        u4_srl_453_n54), .B2(u4_srl_453_n137), .ZN(u4_srl_453_n795) );
  AOI221_X1 u4_srl_453_U796 ( .B1(n6425), .B2(u4_srl_453_n35), .C1(n6422), 
        .C2(u4_srl_453_n41), .A(u4_srl_453_n795), .ZN(u4_srl_453_n571) );
  OAI22_X1 u4_srl_453_U795 ( .A1(u4_srl_453_n653), .A2(u4_srl_453_n168), .B1(
        u4_srl_453_n571), .B2(u4_srl_453_n170), .ZN(u4_srl_453_n793) );
  AOI221_X1 u4_srl_453_U794 ( .B1(u4_srl_453_n162), .B2(u4_srl_453_n253), .C1(
        u4_srl_453_n164), .C2(u4_srl_453_n257), .A(u4_srl_453_n793), .ZN(
        u4_srl_453_n792) );
  AOI21_X1 u4_srl_453_U793 ( .B1(u4_srl_453_n791), .B2(u4_srl_453_n792), .A(
        u4_shift_right[8]), .ZN(u4_N5916) );
  AOI22_X1 u4_srl_453_U792 ( .A1(n6440), .A2(u4_srl_453_n44), .B1(n6431), .B2(
        u4_srl_453_n47), .ZN(u4_srl_453_n790) );
  OAI221_X1 u4_srl_453_U791 ( .B1(u4_srl_453_n31), .B2(u4_srl_453_n144), .C1(
        u4_srl_453_n39), .C2(u4_srl_453_n146), .A(u4_srl_453_n790), .ZN(
        u4_srl_453_n543) );
  AOI22_X1 u4_srl_453_U790 ( .A1(n6429), .A2(u4_srl_453_n44), .B1(n6428), .B2(
        u4_srl_453_n47), .ZN(u4_srl_453_n789) );
  OAI221_X1 u4_srl_453_U789 ( .B1(u4_srl_453_n31), .B2(u4_srl_453_n141), .C1(
        u4_srl_453_n39), .C2(u4_srl_453_n140), .A(u4_srl_453_n789), .ZN(
        u4_srl_453_n638) );
  AOI22_X1 u4_srl_453_U788 ( .A1(n6445), .A2(u4_srl_453_n43), .B1(n6438), .B2(
        u4_srl_453_n47), .ZN(u4_srl_453_n788) );
  OAI221_X1 u4_srl_453_U787 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n151), .C1(
        u4_srl_453_n39), .C2(u4_srl_453_n153), .A(u4_srl_453_n788), .ZN(
        u4_srl_453_n545) );
  AOI22_X1 u4_srl_453_U786 ( .A1(n6436), .A2(u4_srl_453_n45), .B1(n6435), .B2(
        u4_srl_453_n47), .ZN(u4_srl_453_n787) );
  OAI221_X1 u4_srl_453_U785 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n148), .C1(
        u4_srl_453_n38), .C2(u4_srl_453_n147), .A(u4_srl_453_n787), .ZN(
        u4_srl_453_n542) );
  AOI22_X1 u4_srl_453_U784 ( .A1(u4_srl_453_n22), .A2(u4_srl_453_n545), .B1(
        u4_srl_453_n28), .B2(u4_srl_453_n542), .ZN(u4_srl_453_n786) );
  INV_X1 u4_srl_453_U783 ( .A(u4_srl_453_n786), .ZN(u4_srl_453_n785) );
  AOI221_X1 u4_srl_453_U782 ( .B1(u4_srl_453_n543), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n638), .C2(u4_srl_453_n57), .A(u4_srl_453_n785), .ZN(
        u4_srl_453_n449) );
  INV_X1 u4_srl_453_U781 ( .A(u4_srl_453_n449), .ZN(u4_srl_453_n761) );
  AOI22_X1 u4_srl_453_U780 ( .A1(fract_denorm[98]), .A2(u4_srl_453_n44), .B1(
        fract_denorm[97]), .B2(u4_srl_453_n52), .ZN(u4_srl_453_n784) );
  OAI221_X1 u4_srl_453_U779 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n71), .C1(
        u4_srl_453_n38), .C2(u4_srl_453_n73), .A(u4_srl_453_n784), .ZN(
        u4_srl_453_n532) );
  AOI22_X1 u4_srl_453_U778 ( .A1(fract_denorm[94]), .A2(u4_srl_453_n45), .B1(
        fract_denorm[93]), .B2(u4_srl_453_n48), .ZN(u4_srl_453_n783) );
  OAI221_X1 u4_srl_453_U777 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n68), .C1(
        u4_srl_453_n38), .C2(u4_srl_453_n67), .A(u4_srl_453_n783), .ZN(
        u4_srl_453_n527) );
  INV_X1 u4_srl_453_U776 ( .A(u4_srl_453_n247), .ZN(u4_srl_453_n403) );
  AOI22_X1 u4_srl_453_U775 ( .A1(fract_denorm[102]), .A2(u4_srl_453_n44), .B1(
        fract_denorm[101]), .B2(u4_srl_453_n51), .ZN(u4_srl_453_n782) );
  OAI221_X1 u4_srl_453_U774 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n78), .C1(
        u4_srl_453_n38), .C2(u4_srl_453_n75), .A(u4_srl_453_n782), .ZN(
        u4_srl_453_n531) );
  AOI22_X1 u4_srl_453_U773 ( .A1(u4_srl_453_n22), .A2(u4_srl_453_n403), .B1(
        u4_srl_453_n28), .B2(u4_srl_453_n531), .ZN(u4_srl_453_n781) );
  INV_X1 u4_srl_453_U772 ( .A(u4_srl_453_n781), .ZN(u4_srl_453_n780) );
  AOI221_X1 u4_srl_453_U771 ( .B1(u4_srl_453_n532), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n527), .C2(u4_srl_453_n57), .A(u4_srl_453_n780), .ZN(
        u4_srl_453_n189) );
  AOI22_X1 u4_srl_453_U770 ( .A1(fract_denorm[82]), .A2(u4_srl_453_n45), .B1(
        fract_denorm[81]), .B2(u4_srl_453_n47), .ZN(u4_srl_453_n779) );
  OAI221_X1 u4_srl_453_U769 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n97), .C1(
        u4_srl_453_n38), .C2(u4_srl_453_n99), .A(u4_srl_453_n779), .ZN(
        u4_srl_453_n526) );
  INV_X1 u4_srl_453_U768 ( .A(u4_srl_453_n526), .ZN(u4_srl_453_n685) );
  AOI22_X1 u4_srl_453_U767 ( .A1(fract_denorm[78]), .A2(u4_srl_453_n45), .B1(
        fract_denorm[77]), .B2(u4_srl_453_n51), .ZN(u4_srl_453_n778) );
  OAI221_X1 u4_srl_453_U766 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n94), .C1(
        u4_srl_453_n38), .C2(u4_srl_453_n93), .A(u4_srl_453_n778), .ZN(
        u4_srl_453_n628) );
  INV_X1 u4_srl_453_U765 ( .A(u4_srl_453_n628), .ZN(u4_srl_453_n522) );
  AOI22_X1 u4_srl_453_U764 ( .A1(fract_denorm[90]), .A2(u4_srl_453_n45), .B1(
        fract_denorm[89]), .B2(u4_srl_453_n49), .ZN(u4_srl_453_n777) );
  OAI221_X1 u4_srl_453_U763 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n90), .C1(
        u4_srl_453_n38), .C2(u4_srl_453_n92), .A(u4_srl_453_n777), .ZN(
        u4_srl_453_n528) );
  AOI22_X1 u4_srl_453_U762 ( .A1(fract_denorm[86]), .A2(u4_srl_453_n43), .B1(
        fract_denorm[85]), .B2(u4_srl_453_n47), .ZN(u4_srl_453_n776) );
  OAI221_X1 u4_srl_453_U761 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n87), .C1(
        u4_srl_453_n38), .C2(u4_srl_453_n86), .A(u4_srl_453_n776), .ZN(
        u4_srl_453_n525) );
  AOI22_X1 u4_srl_453_U760 ( .A1(u4_srl_453_n22), .A2(u4_srl_453_n528), .B1(
        u4_srl_453_n28), .B2(u4_srl_453_n525), .ZN(u4_srl_453_n775) );
  OAI221_X1 u4_srl_453_U759 ( .B1(u4_srl_453_n685), .B2(u4_srl_453_n19), .C1(
        u4_srl_453_n522), .C2(u4_srl_453_n59), .A(u4_srl_453_n775), .ZN(
        u4_srl_453_n366) );
  INV_X1 u4_srl_453_U758 ( .A(u4_srl_453_n366), .ZN(u4_srl_453_n295) );
  OAI22_X1 u4_srl_453_U757 ( .A1(u4_srl_453_n189), .A2(u4_srl_453_n242), .B1(
        u4_srl_453_n295), .B2(u4_srl_453_n238), .ZN(u4_srl_453_n235) );
  AOI22_X1 u4_srl_453_U756 ( .A1(fract_denorm[66]), .A2(u4_srl_453_n45), .B1(
        fract_denorm[65]), .B2(u4_srl_453_n49), .ZN(u4_srl_453_n774) );
  OAI221_X1 u4_srl_453_U755 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n104), .C1(
        u4_srl_453_n38), .C2(u4_srl_453_n106), .A(u4_srl_453_n774), .ZN(
        u4_srl_453_n538) );
  AOI22_X1 u4_srl_453_U754 ( .A1(fract_denorm[62]), .A2(u4_srl_453_n42), .B1(
        fract_denorm[61]), .B2(u4_srl_453_n47), .ZN(u4_srl_453_n773) );
  OAI221_X1 u4_srl_453_U753 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n101), .C1(
        u4_srl_453_n38), .C2(u4_srl_453_n100), .A(u4_srl_453_n773), .ZN(
        u4_srl_453_n533) );
  AOI22_X1 u4_srl_453_U752 ( .A1(fract_denorm[74]), .A2(u4_srl_453_n43), .B1(
        fract_denorm[73]), .B2(u4_srl_453_n47), .ZN(u4_srl_453_n772) );
  OAI221_X1 u4_srl_453_U751 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n111), .C1(
        u4_srl_453_n38), .C2(u4_srl_453_n113), .A(u4_srl_453_n772), .ZN(
        u4_srl_453_n629) );
  AOI22_X1 u4_srl_453_U750 ( .A1(fract_denorm[70]), .A2(u4_srl_453_n43), .B1(
        fract_denorm[69]), .B2(u4_srl_453_n49), .ZN(u4_srl_453_n771) );
  OAI221_X1 u4_srl_453_U749 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n108), .C1(
        u4_srl_453_n37), .C2(u4_srl_453_n107), .A(u4_srl_453_n771), .ZN(
        u4_srl_453_n537) );
  AOI22_X1 u4_srl_453_U748 ( .A1(u4_srl_453_n22), .A2(u4_srl_453_n629), .B1(
        u4_srl_453_n28), .B2(u4_srl_453_n537), .ZN(u4_srl_453_n770) );
  INV_X1 u4_srl_453_U747 ( .A(u4_srl_453_n770), .ZN(u4_srl_453_n769) );
  AOI221_X1 u4_srl_453_U746 ( .B1(u4_srl_453_n538), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n533), .C2(u4_srl_453_n57), .A(u4_srl_453_n769), .ZN(
        u4_srl_453_n296) );
  AOI22_X1 u4_srl_453_U745 ( .A1(fract_denorm[50]), .A2(u4_srl_453_n43), .B1(
        n6367), .B2(u4_srl_453_n49), .ZN(u4_srl_453_n768) );
  OAI221_X1 u4_srl_453_U744 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n125), .C1(
        u4_srl_453_n37), .C2(u4_srl_453_n126), .A(u4_srl_453_n768), .ZN(
        u4_srl_453_n549) );
  AOI22_X1 u4_srl_453_U743 ( .A1(n6408), .A2(u4_srl_453_n43), .B1(n6407), .B2(
        u4_srl_453_n49), .ZN(u4_srl_453_n767) );
  OAI221_X1 u4_srl_453_U742 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n122), .C1(
        u4_srl_453_n37), .C2(u4_srl_453_n121), .A(u4_srl_453_n767), .ZN(
        u4_srl_453_n544) );
  AOI22_X1 u4_srl_453_U741 ( .A1(fract_denorm[58]), .A2(u4_srl_453_n43), .B1(
        fract_denorm[57]), .B2(u4_srl_453_n49), .ZN(u4_srl_453_n766) );
  OAI221_X1 u4_srl_453_U740 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n83), .C1(
        u4_srl_453_n37), .C2(u4_srl_453_n85), .A(u4_srl_453_n766), .ZN(
        u4_srl_453_n534) );
  AOI22_X1 u4_srl_453_U739 ( .A1(fract_denorm[54]), .A2(u4_srl_453_n43), .B1(
        fract_denorm[53]), .B2(u4_srl_453_n49), .ZN(u4_srl_453_n765) );
  OAI221_X1 u4_srl_453_U738 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n114), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n119), .A(u4_srl_453_n765), .ZN(
        u4_srl_453_n548) );
  AOI22_X1 u4_srl_453_U737 ( .A1(u4_srl_453_n22), .A2(u4_srl_453_n534), .B1(
        u4_srl_453_n28), .B2(u4_srl_453_n548), .ZN(u4_srl_453_n764) );
  INV_X1 u4_srl_453_U736 ( .A(u4_srl_453_n764), .ZN(u4_srl_453_n763) );
  AOI221_X1 u4_srl_453_U735 ( .B1(u4_srl_453_n549), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n544), .C2(u4_srl_453_n57), .A(u4_srl_453_n763), .ZN(
        u4_srl_453_n368) );
  OAI22_X1 u4_srl_453_U734 ( .A1(u4_srl_453_n296), .A2(u4_srl_453_n177), .B1(
        u4_srl_453_n368), .B2(u4_srl_453_n179), .ZN(u4_srl_453_n762) );
  AOI221_X1 u4_srl_453_U733 ( .B1(u4_srl_453_n171), .B2(u4_srl_453_n761), .C1(
        u4_srl_453_n235), .C2(u4_srl_453_n174), .A(u4_srl_453_n762), .ZN(
        u4_srl_453_n754) );
  AOI22_X1 u4_srl_453_U732 ( .A1(n6442), .A2(u4_srl_453_n43), .B1(n6417), .B2(
        u4_srl_453_n49), .ZN(u4_srl_453_n760) );
  OAI221_X1 u4_srl_453_U731 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n131), .C1(
        u4_srl_453_n39), .C2(u4_srl_453_n133), .A(u4_srl_453_n760), .ZN(
        u4_srl_453_n221) );
  AOI22_X1 u4_srl_453_U730 ( .A1(n6415), .A2(u4_srl_453_n43), .B1(n6414), .B2(
        u4_srl_453_n49), .ZN(u4_srl_453_n759) );
  OAI221_X1 u4_srl_453_U729 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n128), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n127), .A(u4_srl_453_n759), .ZN(
        u4_srl_453_n225) );
  OAI22_X1 u4_srl_453_U728 ( .A1(u4_srl_453_n136), .A2(u4_srl_453_n1), .B1(
        u4_srl_453_n135), .B2(u4_srl_453_n54), .ZN(u4_srl_453_n758) );
  AOI221_X1 u4_srl_453_U727 ( .B1(u4_srl_453_n35), .B2(n6420), .C1(
        u4_srl_453_n41), .C2(n6419), .A(u4_srl_453_n758), .ZN(u4_srl_453_n636)
         );
  OAI22_X1 u4_srl_453_U726 ( .A1(u4_srl_453_n155), .A2(u4_srl_453_n1), .B1(
        u4_srl_453_n138), .B2(u4_srl_453_n54), .ZN(u4_srl_453_n757) );
  AOI221_X1 u4_srl_453_U725 ( .B1(n6423), .B2(u4_srl_453_n35), .C1(n6425), 
        .C2(u4_srl_453_n41), .A(u4_srl_453_n757), .ZN(u4_srl_453_n540) );
  OAI22_X1 u4_srl_453_U724 ( .A1(u4_srl_453_n636), .A2(u4_srl_453_n168), .B1(
        u4_srl_453_n540), .B2(u4_srl_453_n170), .ZN(u4_srl_453_n756) );
  AOI221_X1 u4_srl_453_U723 ( .B1(u4_srl_453_n162), .B2(u4_srl_453_n221), .C1(
        u4_srl_453_n164), .C2(u4_srl_453_n225), .A(u4_srl_453_n756), .ZN(
        u4_srl_453_n755) );
  AOI21_X1 u4_srl_453_U722 ( .B1(u4_srl_453_n754), .B2(u4_srl_453_n755), .A(
        u4_shift_right[8]), .ZN(u4_N5917) );
  AOI22_X1 u4_srl_453_U721 ( .A1(u4_srl_453_n22), .A2(u4_srl_453_n514), .B1(
        u4_srl_453_n28), .B2(u4_srl_453_n510), .ZN(u4_srl_453_n753) );
  INV_X1 u4_srl_453_U720 ( .A(u4_srl_453_n753), .ZN(u4_srl_453_n752) );
  AOI221_X1 u4_srl_453_U719 ( .B1(u4_srl_453_n511), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n512), .C2(u4_srl_453_n57), .A(u4_srl_453_n752), .ZN(
        u4_srl_453_n446) );
  INV_X1 u4_srl_453_U718 ( .A(u4_srl_453_n446), .ZN(u4_srl_453_n742) );
  INV_X1 u4_srl_453_U717 ( .A(u4_srl_453_n500), .ZN(u4_srl_453_n750) );
  INV_X1 u4_srl_453_U716 ( .A(u4_srl_453_n605), .ZN(u4_srl_453_n496) );
  AOI22_X1 u4_srl_453_U715 ( .A1(u4_srl_453_n22), .A2(u4_srl_453_n380), .B1(
        u4_srl_453_n28), .B2(u4_srl_453_n499), .ZN(u4_srl_453_n751) );
  OAI221_X1 u4_srl_453_U714 ( .B1(u4_srl_453_n750), .B2(u4_srl_453_n19), .C1(
        u4_srl_453_n496), .C2(u4_srl_453_n59), .A(u4_srl_453_n751), .ZN(
        u4_srl_453_n360) );
  INV_X1 u4_srl_453_U713 ( .A(u4_srl_453_n360), .ZN(u4_srl_453_n188) );
  INV_X1 u4_srl_453_U712 ( .A(u4_srl_453_n601), .ZN(u4_srl_453_n491) );
  AOI22_X1 u4_srl_453_U711 ( .A1(u4_srl_453_n22), .A2(u4_srl_453_n606), .B1(
        u4_srl_453_n28), .B2(u4_srl_453_n494), .ZN(u4_srl_453_n749) );
  OAI221_X1 u4_srl_453_U710 ( .B1(u4_srl_453_n748), .B2(u4_srl_453_n19), .C1(
        u4_srl_453_n491), .C2(u4_srl_453_n59), .A(u4_srl_453_n749), .ZN(
        u4_srl_453_n361) );
  INV_X1 u4_srl_453_U709 ( .A(u4_srl_453_n361), .ZN(u4_srl_453_n279) );
  OAI22_X1 u4_srl_453_U708 ( .A1(u4_srl_453_n188), .A2(u4_srl_453_n242), .B1(
        u4_srl_453_n279), .B2(u4_srl_453_n238), .ZN(u4_srl_453_n234) );
  INV_X1 u4_srl_453_U707 ( .A(u4_srl_453_n609), .ZN(u4_srl_453_n501) );
  AOI22_X1 u4_srl_453_U706 ( .A1(u4_srl_453_n22), .A2(u4_srl_453_n602), .B1(
        u4_srl_453_n28), .B2(u4_srl_453_n504), .ZN(u4_srl_453_n747) );
  OAI221_X1 u4_srl_453_U705 ( .B1(u4_srl_453_n746), .B2(u4_srl_453_n19), .C1(
        u4_srl_453_n501), .C2(u4_srl_453_n59), .A(u4_srl_453_n747), .ZN(
        u4_srl_453_n448) );
  INV_X1 u4_srl_453_U704 ( .A(u4_srl_453_n448), .ZN(u4_srl_453_n280) );
  AOI22_X1 u4_srl_453_U703 ( .A1(u4_srl_453_n22), .A2(u4_srl_453_n506), .B1(
        u4_srl_453_n28), .B2(u4_srl_453_n517), .ZN(u4_srl_453_n745) );
  INV_X1 u4_srl_453_U702 ( .A(u4_srl_453_n745), .ZN(u4_srl_453_n744) );
  AOI221_X1 u4_srl_453_U701 ( .B1(u4_srl_453_n518), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n513), .C2(u4_srl_453_n57), .A(u4_srl_453_n744), .ZN(
        u4_srl_453_n363) );
  OAI22_X1 u4_srl_453_U700 ( .A1(u4_srl_453_n280), .A2(u4_srl_453_n177), .B1(
        u4_srl_453_n363), .B2(u4_srl_453_n179), .ZN(u4_srl_453_n743) );
  AOI221_X1 u4_srl_453_U699 ( .B1(u4_srl_453_n171), .B2(u4_srl_453_n742), .C1(
        u4_srl_453_n234), .C2(u4_srl_453_n174), .A(u4_srl_453_n743), .ZN(
        u4_srl_453_n738) );
  INV_X1 u4_srl_453_U698 ( .A(u4_srl_453_n741), .ZN(u4_srl_453_n508) );
  OAI22_X1 u4_srl_453_U697 ( .A1(u4_srl_453_n197), .A2(u4_srl_453_n168), .B1(
        u4_srl_453_n508), .B2(u4_srl_453_n170), .ZN(u4_srl_453_n740) );
  AOI221_X1 u4_srl_453_U696 ( .B1(u4_srl_453_n162), .B2(u4_srl_453_n327), .C1(
        u4_srl_453_n164), .C2(u4_srl_453_n193), .A(u4_srl_453_n740), .ZN(
        u4_srl_453_n739) );
  AOI21_X1 u4_srl_453_U695 ( .B1(u4_srl_453_n738), .B2(u4_srl_453_n739), .A(
        u4_shift_right[8]), .ZN(u4_N5918) );
  AOI22_X1 u4_srl_453_U694 ( .A1(n6434), .A2(u4_srl_453_n43), .B1(n6433), .B2(
        u4_srl_453_n49), .ZN(u4_srl_453_n737) );
  OAI221_X1 u4_srl_453_U693 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n154), .C1(
        u4_srl_453_n37), .C2(u4_srl_453_n145), .A(u4_srl_453_n737), .ZN(
        u4_srl_453_n481) );
  AOI22_X1 u4_srl_453_U692 ( .A1(n6430), .A2(u4_srl_453_n43), .B1(n6432), .B2(
        u4_srl_453_n49), .ZN(u4_srl_453_n736) );
  OAI221_X1 u4_srl_453_U691 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n143), .C1(
        u4_srl_453_n37), .C2(u4_srl_453_n142), .A(u4_srl_453_n736), .ZN(
        u4_srl_453_n482) );
  AOI22_X1 u4_srl_453_U690 ( .A1(n6406), .A2(u4_srl_453_n43), .B1(n6405), .B2(
        u4_srl_453_n49), .ZN(u4_srl_453_n735) );
  OAI221_X1 u4_srl_453_U689 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n159), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n152), .A(u4_srl_453_n735), .ZN(
        u4_srl_453_n484) );
  AOI22_X1 u4_srl_453_U688 ( .A1(n6437), .A2(u4_srl_453_n43), .B1(n6439), .B2(
        u4_srl_453_n49), .ZN(u4_srl_453_n734) );
  OAI221_X1 u4_srl_453_U687 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n150), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n149), .A(u4_srl_453_n734), .ZN(
        u4_srl_453_n480) );
  AOI22_X1 u4_srl_453_U686 ( .A1(u4_srl_453_n22), .A2(u4_srl_453_n484), .B1(
        u4_srl_453_n27), .B2(u4_srl_453_n480), .ZN(u4_srl_453_n733) );
  INV_X1 u4_srl_453_U685 ( .A(u4_srl_453_n733), .ZN(u4_srl_453_n732) );
  AOI221_X1 u4_srl_453_U684 ( .B1(u4_srl_453_n481), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n482), .C2(u4_srl_453_n57), .A(u4_srl_453_n732), .ZN(
        u4_srl_453_n443) );
  INV_X1 u4_srl_453_U683 ( .A(u4_srl_453_n443), .ZN(u4_srl_453_n709) );
  AOI22_X1 u4_srl_453_U682 ( .A1(fract_denorm[96]), .A2(u4_srl_453_n42), .B1(
        fract_denorm[95]), .B2(u4_srl_453_n49), .ZN(u4_srl_453_n731) );
  OAI221_X1 u4_srl_453_U681 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n70), .C1(
        u4_srl_453_n37), .C2(u4_srl_453_n69), .A(u4_srl_453_n731), .ZN(
        u4_srl_453_n465) );
  AOI22_X1 u4_srl_453_U680 ( .A1(fract_denorm[100]), .A2(u4_srl_453_n45), .B1(
        fract_denorm[99]), .B2(u4_srl_453_n48), .ZN(u4_srl_453_n730) );
  OAI221_X1 u4_srl_453_U679 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n79), .C1(
        u4_srl_453_n37), .C2(u4_srl_453_n72), .A(u4_srl_453_n730), .ZN(
        u4_srl_453_n470) );
  AOI222_X1 u4_srl_453_U678 ( .A1(u4_srl_453_n465), .A2(u4_srl_453_n56), .B1(
        u4_srl_453_n470), .B2(u4_srl_453_n16), .C1(u4_srl_453_n728), .C2(
        u4_srl_453_n729), .ZN(u4_srl_453_n187) );
  AOI22_X1 u4_srl_453_U677 ( .A1(fract_denorm[84]), .A2(u4_srl_453_n45), .B1(
        fract_denorm[83]), .B2(u4_srl_453_n48), .ZN(u4_srl_453_n727) );
  OAI221_X1 u4_srl_453_U676 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n117), .C1(
        u4_srl_453_n37), .C2(u4_srl_453_n98), .A(u4_srl_453_n727), .ZN(
        u4_srl_453_n463) );
  INV_X1 u4_srl_453_U675 ( .A(u4_srl_453_n463), .ZN(u4_srl_453_n663) );
  AOI22_X1 u4_srl_453_U674 ( .A1(fract_denorm[80]), .A2(u4_srl_453_n45), .B1(
        fract_denorm[79]), .B2(u4_srl_453_n48), .ZN(u4_srl_453_n726) );
  OAI221_X1 u4_srl_453_U673 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n96), .C1(
        u4_srl_453_n37), .C2(u4_srl_453_n95), .A(u4_srl_453_n726), .ZN(
        u4_srl_453_n587) );
  INV_X1 u4_srl_453_U672 ( .A(u4_srl_453_n587), .ZN(u4_srl_453_n459) );
  AOI22_X1 u4_srl_453_U671 ( .A1(fract_denorm[92]), .A2(u4_srl_453_n45), .B1(
        fract_denorm[91]), .B2(u4_srl_453_n48), .ZN(u4_srl_453_n725) );
  OAI221_X1 u4_srl_453_U670 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n74), .C1(
        u4_srl_453_n37), .C2(u4_srl_453_n91), .A(u4_srl_453_n725), .ZN(
        u4_srl_453_n466) );
  AOI22_X1 u4_srl_453_U669 ( .A1(fract_denorm[88]), .A2(u4_srl_453_n45), .B1(
        fract_denorm[87]), .B2(u4_srl_453_n48), .ZN(u4_srl_453_n724) );
  OAI221_X1 u4_srl_453_U668 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n89), .C1(
        u4_srl_453_n37), .C2(u4_srl_453_n88), .A(u4_srl_453_n724), .ZN(
        u4_srl_453_n462) );
  AOI22_X1 u4_srl_453_U667 ( .A1(u4_srl_453_n22), .A2(u4_srl_453_n466), .B1(
        u4_srl_453_n27), .B2(u4_srl_453_n462), .ZN(u4_srl_453_n723) );
  OAI221_X1 u4_srl_453_U666 ( .B1(u4_srl_453_n663), .B2(u4_srl_453_n19), .C1(
        u4_srl_453_n459), .C2(u4_srl_453_n59), .A(u4_srl_453_n723), .ZN(
        u4_srl_453_n356) );
  INV_X1 u4_srl_453_U665 ( .A(u4_srl_453_n356), .ZN(u4_srl_453_n277) );
  OAI22_X1 u4_srl_453_U664 ( .A1(u4_srl_453_n187), .A2(u4_srl_453_n242), .B1(
        u4_srl_453_n277), .B2(u4_srl_453_n238), .ZN(u4_srl_453_n233) );
  AOI22_X1 u4_srl_453_U663 ( .A1(fract_denorm[68]), .A2(u4_srl_453_n45), .B1(
        fract_denorm[67]), .B2(u4_srl_453_n48), .ZN(u4_srl_453_n722) );
  OAI221_X1 u4_srl_453_U662 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n116), .C1(
        u4_srl_453_n37), .C2(u4_srl_453_n105), .A(u4_srl_453_n722), .ZN(
        u4_srl_453_n476) );
  AOI22_X1 u4_srl_453_U661 ( .A1(fract_denorm[64]), .A2(u4_srl_453_n45), .B1(
        fract_denorm[63]), .B2(u4_srl_453_n48), .ZN(u4_srl_453_n721) );
  OAI221_X1 u4_srl_453_U660 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n103), .C1(
        u4_srl_453_n37), .C2(u4_srl_453_n102), .A(u4_srl_453_n721), .ZN(
        u4_srl_453_n471) );
  AOI22_X1 u4_srl_453_U659 ( .A1(fract_denorm[76]), .A2(u4_srl_453_n42), .B1(
        fract_denorm[75]), .B2(u4_srl_453_n48), .ZN(u4_srl_453_n720) );
  OAI221_X1 u4_srl_453_U658 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n118), .C1(
        u4_srl_453_n37), .C2(u4_srl_453_n112), .A(u4_srl_453_n720), .ZN(
        u4_srl_453_n588) );
  AOI22_X1 u4_srl_453_U657 ( .A1(fract_denorm[72]), .A2(u4_srl_453_n45), .B1(
        fract_denorm[71]), .B2(u4_srl_453_n48), .ZN(u4_srl_453_n719) );
  OAI221_X1 u4_srl_453_U656 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n110), .C1(
        u4_srl_453_n37), .C2(u4_srl_453_n109), .A(u4_srl_453_n719), .ZN(
        u4_srl_453_n475) );
  AOI22_X1 u4_srl_453_U655 ( .A1(u4_srl_453_n20), .A2(u4_srl_453_n588), .B1(
        u4_srl_453_n27), .B2(u4_srl_453_n475), .ZN(u4_srl_453_n718) );
  INV_X1 u4_srl_453_U654 ( .A(u4_srl_453_n718), .ZN(u4_srl_453_n717) );
  AOI221_X1 u4_srl_453_U653 ( .B1(u4_srl_453_n476), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n471), .C2(u4_srl_453_n57), .A(u4_srl_453_n717), .ZN(
        u4_srl_453_n278) );
  AOI22_X1 u4_srl_453_U652 ( .A1(fract_denorm[52]), .A2(u4_srl_453_n45), .B1(
        fract_denorm[51]), .B2(u4_srl_453_n48), .ZN(u4_srl_453_n716) );
  OAI221_X1 u4_srl_453_U651 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n120), .C1(
        u4_srl_453_n37), .C2(u4_srl_453_n80), .A(u4_srl_453_n716), .ZN(
        u4_srl_453_n488) );
  AOI22_X1 u4_srl_453_U650 ( .A1(n6409), .A2(u4_srl_453_n45), .B1(n6410), .B2(
        u4_srl_453_n48), .ZN(u4_srl_453_n715) );
  OAI221_X1 u4_srl_453_U649 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n124), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n123), .A(u4_srl_453_n715), .ZN(
        u4_srl_453_n483) );
  AOI22_X1 u4_srl_453_U648 ( .A1(fract_denorm[60]), .A2(u4_srl_453_n42), .B1(
        fract_denorm[59]), .B2(u4_srl_453_n48), .ZN(u4_srl_453_n714) );
  OAI221_X1 u4_srl_453_U647 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n115), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n84), .A(u4_srl_453_n714), .ZN(
        u4_srl_453_n472) );
  AOI22_X1 u4_srl_453_U646 ( .A1(fract_denorm[56]), .A2(u4_srl_453_n42), .B1(
        fract_denorm[55]), .B2(u4_srl_453_n47), .ZN(u4_srl_453_n713) );
  OAI221_X1 u4_srl_453_U645 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n82), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n81), .A(u4_srl_453_n713), .ZN(
        u4_srl_453_n487) );
  AOI22_X1 u4_srl_453_U644 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n472), .B1(
        u4_srl_453_n27), .B2(u4_srl_453_n487), .ZN(u4_srl_453_n712) );
  INV_X1 u4_srl_453_U643 ( .A(u4_srl_453_n712), .ZN(u4_srl_453_n711) );
  AOI221_X1 u4_srl_453_U642 ( .B1(u4_srl_453_n488), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n483), .C2(u4_srl_453_n57), .A(u4_srl_453_n711), .ZN(
        u4_srl_453_n358) );
  OAI22_X1 u4_srl_453_U641 ( .A1(u4_srl_453_n278), .A2(u4_srl_453_n177), .B1(
        u4_srl_453_n358), .B2(u4_srl_453_n179), .ZN(u4_srl_453_n710) );
  AOI221_X1 u4_srl_453_U640 ( .B1(u4_srl_453_n171), .B2(u4_srl_453_n709), .C1(
        u4_srl_453_n233), .C2(u4_srl_453_n174), .A(u4_srl_453_n710), .ZN(
        u4_srl_453_n702) );
  AOI22_X1 u4_srl_453_U639 ( .A1(n6420), .A2(u4_srl_453_n42), .B1(n6419), .B2(
        u4_srl_453_n47), .ZN(u4_srl_453_n708) );
  OAI221_X1 u4_srl_453_U638 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n156), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n132), .A(u4_srl_453_n708), .ZN(
        u4_srl_453_n283) );
  AOI22_X1 u4_srl_453_U637 ( .A1(n6416), .A2(u4_srl_453_n42), .B1(n6418), .B2(
        u4_srl_453_n47), .ZN(u4_srl_453_n707) );
  OAI221_X1 u4_srl_453_U636 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n130), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n129), .A(u4_srl_453_n707), .ZN(
        u4_srl_453_n163) );
  OAI22_X1 u4_srl_453_U635 ( .A1(u4_srl_453_n137), .A2(u4_srl_453_n1), .B1(
        u4_srl_453_n139), .B2(u4_srl_453_n54), .ZN(u4_srl_453_n706) );
  AOI221_X1 u4_srl_453_U634 ( .B1(u4_srl_453_n35), .B2(n6422), .C1(
        u4_srl_453_n41), .C2(n6421), .A(u4_srl_453_n706), .ZN(u4_srl_453_n169)
         );
  AOI22_X1 u4_srl_453_U633 ( .A1(n6427), .A2(u4_srl_453_n42), .B1(n6426), .B2(
        u4_srl_453_n47), .ZN(u4_srl_453_n705) );
  OAI221_X1 u4_srl_453_U632 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n155), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n138), .A(u4_srl_453_n705), .ZN(
        u4_srl_453_n670) );
  INV_X1 u4_srl_453_U631 ( .A(u4_srl_453_n670), .ZN(u4_srl_453_n478) );
  OAI22_X1 u4_srl_453_U630 ( .A1(u4_srl_453_n169), .A2(u4_srl_453_n168), .B1(
        u4_srl_453_n478), .B2(u4_srl_453_n170), .ZN(u4_srl_453_n704) );
  AOI221_X1 u4_srl_453_U629 ( .B1(u4_srl_453_n162), .B2(u4_srl_453_n283), .C1(
        u4_srl_453_n164), .C2(u4_srl_453_n163), .A(u4_srl_453_n704), .ZN(
        u4_srl_453_n703) );
  AOI21_X1 u4_srl_453_U628 ( .B1(u4_srl_453_n702), .B2(u4_srl_453_n703), .A(
        u4_shift_right[8]), .ZN(u4_N5919) );
  AOI22_X1 u4_srl_453_U627 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n575), .B1(
        u4_srl_453_n27), .B2(u4_srl_453_n576), .ZN(u4_srl_453_n701) );
  INV_X1 u4_srl_453_U626 ( .A(u4_srl_453_n701), .ZN(u4_srl_453_n700) );
  AOI221_X1 u4_srl_453_U625 ( .B1(u4_srl_453_n573), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n574), .C2(u4_srl_453_n57), .A(u4_srl_453_n700), .ZN(
        u4_srl_453_n429) );
  INV_X1 u4_srl_453_U624 ( .A(u4_srl_453_n429), .ZN(u4_srl_453_n692) );
  AOI222_X1 u4_srl_453_U623 ( .A1(u4_srl_453_n562), .A2(u4_srl_453_n15), .B1(
        u4_srl_453_n406), .B2(u4_srl_453_n25), .C1(u4_srl_453_n563), .C2(
        u4_srl_453_n56), .ZN(u4_srl_453_n186) );
  INV_X1 u4_srl_453_U622 ( .A(u4_srl_453_n556), .ZN(u4_srl_453_n648) );
  AOI22_X1 u4_srl_453_U621 ( .A1(u4_srl_453_n20), .A2(u4_srl_453_n558), .B1(
        u4_srl_453_n27), .B2(u4_srl_453_n559), .ZN(u4_srl_453_n699) );
  OAI221_X1 u4_srl_453_U620 ( .B1(u4_srl_453_n648), .B2(u4_srl_453_n19), .C1(
        u4_srl_453_n698), .C2(u4_srl_453_n58), .A(u4_srl_453_n699), .ZN(
        u4_srl_453_n432) );
  INV_X1 u4_srl_453_U619 ( .A(u4_srl_453_n432), .ZN(u4_srl_453_n275) );
  OAI22_X1 u4_srl_453_U618 ( .A1(u4_srl_453_n186), .A2(u4_srl_453_n242), .B1(
        u4_srl_453_n275), .B2(u4_srl_453_n238), .ZN(u4_srl_453_n232) );
  AOI22_X1 u4_srl_453_U617 ( .A1(u4_srl_453_n20), .A2(u4_srl_453_n645), .B1(
        u4_srl_453_n27), .B2(u4_srl_453_n646), .ZN(u4_srl_453_n697) );
  INV_X1 u4_srl_453_U616 ( .A(u4_srl_453_n697), .ZN(u4_srl_453_n696) );
  AOI221_X1 u4_srl_453_U615 ( .B1(u4_srl_453_n568), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n569), .C2(u4_srl_453_n57), .A(u4_srl_453_n696), .ZN(
        u4_srl_453_n276) );
  AOI22_X1 u4_srl_453_U614 ( .A1(u4_srl_453_n20), .A2(u4_srl_453_n564), .B1(
        u4_srl_453_n27), .B2(u4_srl_453_n565), .ZN(u4_srl_453_n695) );
  INV_X1 u4_srl_453_U613 ( .A(u4_srl_453_n695), .ZN(u4_srl_453_n694) );
  AOI221_X1 u4_srl_453_U612 ( .B1(u4_srl_453_n579), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n580), .C2(u4_srl_453_n57), .A(u4_srl_453_n694), .ZN(
        u4_srl_453_n353) );
  OAI22_X1 u4_srl_453_U611 ( .A1(u4_srl_453_n276), .A2(u4_srl_453_n177), .B1(
        u4_srl_453_n353), .B2(u4_srl_453_n179), .ZN(u4_srl_453_n693) );
  AOI221_X1 u4_srl_453_U610 ( .B1(u4_srl_453_n171), .B2(u4_srl_453_n692), .C1(
        u4_srl_453_n232), .C2(u4_srl_453_n174), .A(u4_srl_453_n693), .ZN(
        u4_srl_453_n689) );
  INV_X1 u4_srl_453_U609 ( .A(u4_srl_453_n655), .ZN(u4_srl_453_n570) );
  OAI22_X1 u4_srl_453_U608 ( .A1(u4_srl_453_n571), .A2(u4_srl_453_n168), .B1(
        u4_srl_453_n570), .B2(u4_srl_453_n170), .ZN(u4_srl_453_n691) );
  AOI221_X1 u4_srl_453_U607 ( .B1(u4_srl_453_n162), .B2(u4_srl_453_n252), .C1(
        u4_srl_453_n164), .C2(u4_srl_453_n253), .A(u4_srl_453_n691), .ZN(
        u4_srl_453_n690) );
  AOI21_X1 u4_srl_453_U606 ( .B1(u4_srl_453_n689), .B2(u4_srl_453_n690), .A(
        u4_shift_right[8]), .ZN(u4_N5920) );
  AOI22_X1 u4_srl_453_U605 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n544), .B1(
        u4_srl_453_n27), .B2(u4_srl_453_n545), .ZN(u4_srl_453_n688) );
  INV_X1 u4_srl_453_U604 ( .A(u4_srl_453_n688), .ZN(u4_srl_453_n687) );
  AOI221_X1 u4_srl_453_U603 ( .B1(u4_srl_453_n542), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n543), .C2(u4_srl_453_n57), .A(u4_srl_453_n687), .ZN(
        u4_srl_453_n424) );
  INV_X1 u4_srl_453_U602 ( .A(u4_srl_453_n424), .ZN(u4_srl_453_n679) );
  AOI222_X1 u4_srl_453_U601 ( .A1(u4_srl_453_n531), .A2(u4_srl_453_n15), .B1(
        u4_srl_453_n403), .B2(u4_srl_453_n25), .C1(u4_srl_453_n532), .C2(
        u4_srl_453_n56), .ZN(u4_srl_453_n185) );
  INV_X1 u4_srl_453_U600 ( .A(u4_srl_453_n525), .ZN(u4_srl_453_n631) );
  AOI22_X1 u4_srl_453_U599 ( .A1(u4_srl_453_n20), .A2(u4_srl_453_n527), .B1(
        u4_srl_453_n27), .B2(u4_srl_453_n528), .ZN(u4_srl_453_n686) );
  OAI221_X1 u4_srl_453_U598 ( .B1(u4_srl_453_n631), .B2(u4_srl_453_n19), .C1(
        u4_srl_453_n685), .C2(u4_srl_453_n58), .A(u4_srl_453_n686), .ZN(
        u4_srl_453_n427) );
  INV_X1 u4_srl_453_U597 ( .A(u4_srl_453_n427), .ZN(u4_srl_453_n273) );
  OAI22_X1 u4_srl_453_U596 ( .A1(u4_srl_453_n185), .A2(u4_srl_453_n242), .B1(
        u4_srl_453_n273), .B2(u4_srl_453_n238), .ZN(u4_srl_453_n231) );
  INV_X1 u4_srl_453_U595 ( .A(u4_srl_453_n537), .ZN(u4_srl_453_n626) );
  INV_X1 u4_srl_453_U594 ( .A(u4_srl_453_n538), .ZN(u4_srl_453_n683) );
  AOI22_X1 u4_srl_453_U593 ( .A1(u4_srl_453_n20), .A2(u4_srl_453_n628), .B1(
        u4_srl_453_n27), .B2(u4_srl_453_n629), .ZN(u4_srl_453_n684) );
  OAI221_X1 u4_srl_453_U592 ( .B1(u4_srl_453_n626), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n683), .C2(u4_srl_453_n58), .A(u4_srl_453_n684), .ZN(
        u4_srl_453_n426) );
  INV_X1 u4_srl_453_U591 ( .A(u4_srl_453_n426), .ZN(u4_srl_453_n274) );
  AOI22_X1 u4_srl_453_U590 ( .A1(u4_srl_453_n20), .A2(u4_srl_453_n533), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n534), .ZN(u4_srl_453_n682) );
  INV_X1 u4_srl_453_U589 ( .A(u4_srl_453_n682), .ZN(u4_srl_453_n681) );
  AOI221_X1 u4_srl_453_U588 ( .B1(u4_srl_453_n548), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n549), .C2(u4_srl_453_n57), .A(u4_srl_453_n681), .ZN(
        u4_srl_453_n350) );
  OAI22_X1 u4_srl_453_U587 ( .A1(u4_srl_453_n274), .A2(u4_srl_453_n177), .B1(
        u4_srl_453_n350), .B2(u4_srl_453_n179), .ZN(u4_srl_453_n680) );
  AOI221_X1 u4_srl_453_U586 ( .B1(u4_srl_453_n171), .B2(u4_srl_453_n679), .C1(
        u4_srl_453_n231), .C2(u4_srl_453_n174), .A(u4_srl_453_n680), .ZN(
        u4_srl_453_n676) );
  INV_X1 u4_srl_453_U585 ( .A(u4_srl_453_n636), .ZN(u4_srl_453_n219) );
  INV_X1 u4_srl_453_U584 ( .A(u4_srl_453_n638), .ZN(u4_srl_453_n539) );
  OAI22_X1 u4_srl_453_U583 ( .A1(u4_srl_453_n540), .A2(u4_srl_453_n168), .B1(
        u4_srl_453_n539), .B2(u4_srl_453_n170), .ZN(u4_srl_453_n678) );
  AOI221_X1 u4_srl_453_U582 ( .B1(u4_srl_453_n162), .B2(u4_srl_453_n219), .C1(
        u4_srl_453_n164), .C2(u4_srl_453_n221), .A(u4_srl_453_n678), .ZN(
        u4_srl_453_n677) );
  AOI21_X1 u4_srl_453_U581 ( .B1(u4_srl_453_n676), .B2(u4_srl_453_n677), .A(
        u4_shift_right[8]), .ZN(u4_N5921) );
  AOI22_X1 u4_srl_453_U580 ( .A1(u4_srl_453_n346), .A2(u4_srl_453_n401), .B1(
        u4_srl_453_n347), .B2(u4_srl_453_n400), .ZN(u4_srl_453_n215) );
  INV_X1 u4_srl_453_U579 ( .A(u4_srl_453_n423), .ZN(u4_srl_453_n343) );
  OAI222_X1 u4_srl_453_U578 ( .A1(u4_srl_453_n4), .A2(u4_srl_453_n344), .B1(
        u4_srl_453_n383), .B2(u4_srl_453_n215), .C1(u4_srl_453_n11), .C2(
        u4_srl_453_n343), .ZN(u4_srl_453_n675) );
  INV_X1 u4_srl_453_U577 ( .A(u4_srl_453_n675), .ZN(u4_srl_453_n674) );
  OAI221_X1 u4_srl_453_U576 ( .B1(u4_srl_453_n421), .B2(u4_srl_453_n9), .C1(
        u4_srl_453_n673), .C2(u4_srl_453_n8), .A(u4_srl_453_n674), .ZN(
        u4_N5922) );
  AOI22_X1 u4_srl_453_U575 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n483), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n484), .ZN(u4_srl_453_n672) );
  INV_X1 u4_srl_453_U574 ( .A(u4_srl_453_n672), .ZN(u4_srl_453_n671) );
  AOI221_X1 u4_srl_453_U573 ( .B1(u4_srl_453_n480), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n481), .C2(u4_srl_453_n57), .A(u4_srl_453_n671), .ZN(
        u4_srl_453_n418) );
  INV_X1 u4_srl_453_U572 ( .A(u4_srl_453_n283), .ZN(u4_srl_453_n167) );
  AOI22_X1 u4_srl_453_U571 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n482), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n670), .ZN(u4_srl_453_n669) );
  OAI221_X1 u4_srl_453_U570 ( .B1(u4_srl_453_n169), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n167), .C2(u4_srl_453_n58), .A(u4_srl_453_n669), .ZN(
        u4_srl_453_n668) );
  INV_X1 u4_srl_453_U569 ( .A(u4_srl_453_n668), .ZN(u4_srl_453_n618) );
  AOI22_X1 u4_srl_453_U568 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n471), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n472), .ZN(u4_srl_453_n667) );
  INV_X1 u4_srl_453_U567 ( .A(u4_srl_453_n667), .ZN(u4_srl_453_n666) );
  AOI221_X1 u4_srl_453_U566 ( .B1(u4_srl_453_n487), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n488), .C2(u4_srl_453_n57), .A(u4_srl_453_n666), .ZN(
        u4_srl_453_n339) );
  AOI222_X1 u4_srl_453_U565 ( .A1(u4_srl_453_n469), .A2(u4_srl_453_n15), .B1(
        u4_srl_453_n25), .B2(u4_srl_453_n665), .C1(u4_srl_453_n470), .C2(
        u4_srl_453_n56), .ZN(u4_srl_453_n183) );
  INV_X1 u4_srl_453_U564 ( .A(u4_srl_453_n183), .ZN(u4_srl_453_n341) );
  INV_X1 u4_srl_453_U563 ( .A(u4_srl_453_n462), .ZN(u4_srl_453_n662) );
  AOI22_X1 u4_srl_453_U562 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n465), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n466), .ZN(u4_srl_453_n664) );
  OAI221_X1 u4_srl_453_U561 ( .B1(u4_srl_453_n662), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n663), .C2(u4_srl_453_n58), .A(u4_srl_453_n664), .ZN(
        u4_srl_453_n342) );
  AOI22_X1 u4_srl_453_U560 ( .A1(u4_srl_453_n341), .A2(u4_srl_453_n401), .B1(
        u4_srl_453_n342), .B2(u4_srl_453_n400), .ZN(u4_srl_453_n214) );
  AOI22_X1 u4_srl_453_U559 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n587), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n588), .ZN(u4_srl_453_n661) );
  INV_X1 u4_srl_453_U558 ( .A(u4_srl_453_n661), .ZN(u4_srl_453_n660) );
  AOI221_X1 u4_srl_453_U557 ( .B1(u4_srl_453_n475), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n476), .C2(u4_srl_453_n57), .A(u4_srl_453_n660), .ZN(
        u4_srl_453_n338) );
  OAI222_X1 u4_srl_453_U556 ( .A1(u4_srl_453_n4), .A2(u4_srl_453_n339), .B1(
        u4_srl_453_n383), .B2(u4_srl_453_n214), .C1(u4_srl_453_n11), .C2(
        u4_srl_453_n338), .ZN(u4_srl_453_n659) );
  INV_X1 u4_srl_453_U555 ( .A(u4_srl_453_n659), .ZN(u4_srl_453_n658) );
  OAI221_X1 u4_srl_453_U554 ( .B1(u4_srl_453_n418), .B2(u4_srl_453_n10), .C1(
        u4_srl_453_n618), .C2(u4_srl_453_n8), .A(u4_srl_453_n658), .ZN(
        u4_N5923) );
  AOI22_X1 u4_srl_453_U553 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n580), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n575), .ZN(u4_srl_453_n657) );
  INV_X1 u4_srl_453_U552 ( .A(u4_srl_453_n657), .ZN(u4_srl_453_n656) );
  AOI221_X1 u4_srl_453_U551 ( .B1(u4_srl_453_n576), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n573), .C2(u4_srl_453_n57), .A(u4_srl_453_n656), .ZN(
        u4_srl_453_n415) );
  AOI22_X1 u4_srl_453_U550 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n574), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n655), .ZN(u4_srl_453_n654) );
  OAI221_X1 u4_srl_453_U549 ( .B1(u4_srl_453_n571), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n653), .C2(u4_srl_453_n58), .A(u4_srl_453_n654), .ZN(
        u4_srl_453_n652) );
  INV_X1 u4_srl_453_U548 ( .A(u4_srl_453_n652), .ZN(u4_srl_453_n439) );
  AOI22_X1 u4_srl_453_U547 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n569), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n564), .ZN(u4_srl_453_n651) );
  INV_X1 u4_srl_453_U546 ( .A(u4_srl_453_n651), .ZN(u4_srl_453_n650) );
  AOI221_X1 u4_srl_453_U545 ( .B1(u4_srl_453_n565), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n579), .C2(u4_srl_453_n57), .A(u4_srl_453_n650), .ZN(
        u4_srl_453_n321) );
  AOI22_X1 u4_srl_453_U544 ( .A1(u4_srl_453_n562), .A2(u4_srl_453_n409), .B1(
        u4_srl_453_n406), .B2(u4_srl_453_n16), .ZN(u4_srl_453_n182) );
  INV_X1 u4_srl_453_U543 ( .A(u4_srl_453_n182), .ZN(u4_srl_453_n323) );
  INV_X1 u4_srl_453_U542 ( .A(u4_srl_453_n559), .ZN(u4_srl_453_n647) );
  AOI22_X1 u4_srl_453_U541 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n563), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n558), .ZN(u4_srl_453_n649) );
  OAI221_X1 u4_srl_453_U540 ( .B1(u4_srl_453_n647), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n648), .C2(u4_srl_453_n59), .A(u4_srl_453_n649), .ZN(
        u4_srl_453_n324) );
  AOI22_X1 u4_srl_453_U539 ( .A1(u4_srl_453_n323), .A2(u4_srl_453_n401), .B1(
        u4_srl_453_n324), .B2(u4_srl_453_n400), .ZN(u4_srl_453_n213) );
  INV_X1 u4_srl_453_U538 ( .A(u4_srl_453_n646), .ZN(u4_srl_453_n554) );
  INV_X1 u4_srl_453_U537 ( .A(u4_srl_453_n568), .ZN(u4_srl_453_n643) );
  AOI22_X1 u4_srl_453_U536 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n557), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n645), .ZN(u4_srl_453_n644) );
  OAI221_X1 u4_srl_453_U535 ( .B1(u4_srl_453_n554), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n643), .C2(u4_srl_453_n59), .A(u4_srl_453_n644), .ZN(
        u4_srl_453_n417) );
  INV_X1 u4_srl_453_U534 ( .A(u4_srl_453_n417), .ZN(u4_srl_453_n320) );
  OAI222_X1 u4_srl_453_U533 ( .A1(u4_srl_453_n4), .A2(u4_srl_453_n321), .B1(
        u4_srl_453_n383), .B2(u4_srl_453_n213), .C1(u4_srl_453_n11), .C2(
        u4_srl_453_n320), .ZN(u4_srl_453_n642) );
  INV_X1 u4_srl_453_U532 ( .A(u4_srl_453_n642), .ZN(u4_srl_453_n641) );
  OAI221_X1 u4_srl_453_U531 ( .B1(u4_srl_453_n415), .B2(u4_srl_453_n10), .C1(
        u4_srl_453_n439), .C2(u4_srl_453_n8), .A(u4_srl_453_n641), .ZN(
        u4_N5924) );
  AOI22_X1 u4_srl_453_U530 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n549), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n544), .ZN(u4_srl_453_n640) );
  INV_X1 u4_srl_453_U529 ( .A(u4_srl_453_n640), .ZN(u4_srl_453_n639) );
  AOI221_X1 u4_srl_453_U528 ( .B1(u4_srl_453_n545), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n542), .C2(u4_srl_453_n57), .A(u4_srl_453_n639), .ZN(
        u4_srl_453_n398) );
  AOI22_X1 u4_srl_453_U527 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n543), .B1(
        u4_srl_453_n28), .B2(u4_srl_453_n638), .ZN(u4_srl_453_n637) );
  OAI221_X1 u4_srl_453_U526 ( .B1(u4_srl_453_n540), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n636), .C2(u4_srl_453_n59), .A(u4_srl_453_n637), .ZN(
        u4_srl_453_n635) );
  INV_X1 u4_srl_453_U525 ( .A(u4_srl_453_n635), .ZN(u4_srl_453_n390) );
  AOI22_X1 u4_srl_453_U524 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n538), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n533), .ZN(u4_srl_453_n634) );
  INV_X1 u4_srl_453_U523 ( .A(u4_srl_453_n634), .ZN(u4_srl_453_n633) );
  AOI221_X1 u4_srl_453_U522 ( .B1(u4_srl_453_n534), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n548), .C2(u4_srl_453_n57), .A(u4_srl_453_n633), .ZN(
        u4_srl_453_n316) );
  AOI22_X1 u4_srl_453_U521 ( .A1(u4_srl_453_n531), .A2(u4_srl_453_n409), .B1(
        u4_srl_453_n403), .B2(u4_srl_453_n16), .ZN(u4_srl_453_n180) );
  INV_X1 u4_srl_453_U520 ( .A(u4_srl_453_n180), .ZN(u4_srl_453_n318) );
  INV_X1 u4_srl_453_U519 ( .A(u4_srl_453_n528), .ZN(u4_srl_453_n630) );
  AOI22_X1 u4_srl_453_U518 ( .A1(u4_srl_453_n20), .A2(u4_srl_453_n532), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n527), .ZN(u4_srl_453_n632) );
  OAI221_X1 u4_srl_453_U517 ( .B1(u4_srl_453_n630), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n631), .C2(u4_srl_453_n59), .A(u4_srl_453_n632), .ZN(
        u4_srl_453_n319) );
  AOI22_X1 u4_srl_453_U516 ( .A1(u4_srl_453_n318), .A2(u4_srl_453_n401), .B1(
        u4_srl_453_n319), .B2(u4_srl_453_n400), .ZN(u4_srl_453_n211) );
  INV_X1 u4_srl_453_U515 ( .A(u4_srl_453_n629), .ZN(u4_srl_453_n523) );
  AOI22_X1 u4_srl_453_U514 ( .A1(u4_srl_453_n20), .A2(u4_srl_453_n526), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n628), .ZN(u4_srl_453_n627) );
  OAI221_X1 u4_srl_453_U513 ( .B1(u4_srl_453_n523), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n626), .C2(u4_srl_453_n59), .A(u4_srl_453_n627), .ZN(
        u4_srl_453_n399) );
  INV_X1 u4_srl_453_U512 ( .A(u4_srl_453_n399), .ZN(u4_srl_453_n315) );
  OAI222_X1 u4_srl_453_U511 ( .A1(u4_srl_453_n4), .A2(u4_srl_453_n316), .B1(
        u4_srl_453_n383), .B2(u4_srl_453_n211), .C1(u4_srl_453_n11), .C2(
        u4_srl_453_n315), .ZN(u4_srl_453_n625) );
  INV_X1 u4_srl_453_U510 ( .A(u4_srl_453_n625), .ZN(u4_srl_453_n624) );
  OAI221_X1 u4_srl_453_U509 ( .B1(u4_srl_453_n398), .B2(u4_srl_453_n9), .C1(
        u4_srl_453_n390), .C2(u4_srl_453_n8), .A(u4_srl_453_n624), .ZN(
        u4_N5925) );
  INV_X1 u4_srl_453_U508 ( .A(u4_srl_453_n338), .ZN(u4_srl_453_n420) );
  AOI222_X1 u4_srl_453_U507 ( .A1(u4_srl_453_n420), .A2(u4_srl_453_n400), .B1(
        u4_srl_453_n341), .B2(u4_srl_453_n336), .C1(u4_srl_453_n342), .C2(
        u4_srl_453_n401), .ZN(u4_srl_453_n271) );
  INV_X1 u4_srl_453_U506 ( .A(u4_srl_453_n418), .ZN(u4_srl_453_n614) );
  AOI22_X1 u4_srl_453_U505 ( .A1(u4_srl_453_n41), .A2(n6344), .B1(
        u4_srl_453_n35), .B2(n6345), .ZN(u4_srl_453_n623) );
  INV_X1 u4_srl_453_U504 ( .A(u4_srl_453_n623), .ZN(u4_srl_453_n622) );
  AOI221_X1 u4_srl_453_U503 ( .B1(n6347), .B2(u4_srl_453_n42), .C1(n6346), 
        .C2(u4_srl_453_n47), .A(u4_srl_453_n622), .ZN(u4_srl_453_n616) );
  AOI22_X1 u4_srl_453_U502 ( .A1(n6351), .A2(u4_srl_453_n42), .B1(n6350), .B2(
        u4_srl_453_n47), .ZN(u4_srl_453_n621) );
  OAI221_X1 u4_srl_453_U501 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n64), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n63), .A(u4_srl_453_n621), .ZN(
        u4_srl_453_n286) );
  AOI22_X1 u4_srl_453_U500 ( .A1(n6413), .A2(u4_srl_453_n42), .B1(n6411), .B2(
        u4_srl_453_n47), .ZN(u4_srl_453_n620) );
  OAI221_X1 u4_srl_453_U499 ( .B1(u4_srl_453_n30), .B2(u4_srl_453_n157), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n158), .A(u4_srl_453_n620), .ZN(
        u4_srl_453_n165) );
  AOI222_X1 u4_srl_453_U498 ( .A1(u4_srl_453_n15), .A2(u4_srl_453_n286), .B1(
        u4_srl_453_n21), .B2(u4_srl_453_n163), .C1(u4_srl_453_n25), .C2(
        u4_srl_453_n165), .ZN(u4_srl_453_n619) );
  MUX2_X1 u4_srl_453_U497 ( .A(u4_srl_453_n618), .B(u4_srl_453_n619), .S(
        u4_srl_453_n392), .Z(u4_srl_453_n617) );
  OAI21_X1 u4_srl_453_U496 ( .B1(u4_srl_453_n616), .B2(u4_srl_453_n265), .A(
        u4_srl_453_n617), .ZN(u4_srl_453_n615) );
  AOI22_X1 u4_srl_453_U495 ( .A1(u4_srl_453_n14), .A2(u4_srl_453_n614), .B1(
        u4_srl_453_n386), .B2(u4_srl_453_n615), .ZN(u4_srl_453_n613) );
  OAI221_X1 u4_srl_453_U494 ( .B1(u4_srl_453_n271), .B2(u4_srl_453_n383), .C1(
        u4_srl_453_n339), .C2(u4_srl_453_n11), .A(u4_srl_453_n613), .ZN(
        u4_N5907) );
  AOI22_X1 u4_srl_453_U493 ( .A1(u4_srl_453_n20), .A2(u4_srl_453_n518), .B1(
        u4_srl_453_n28), .B2(u4_srl_453_n513), .ZN(u4_srl_453_n612) );
  INV_X1 u4_srl_453_U492 ( .A(u4_srl_453_n612), .ZN(u4_srl_453_n611) );
  AOI221_X1 u4_srl_453_U491 ( .B1(u4_srl_453_n514), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n510), .C2(u4_srl_453_n57), .A(u4_srl_453_n611), .ZN(
        u4_srl_453_n333) );
  AOI22_X1 u4_srl_453_U490 ( .A1(u4_srl_453_n20), .A2(u4_srl_453_n511), .B1(
        u4_srl_453_n28), .B2(u4_srl_453_n512), .ZN(u4_srl_453_n610) );
  OAI221_X1 u4_srl_453_U489 ( .B1(u4_srl_453_n508), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n197), .C2(u4_srl_453_n59), .A(u4_srl_453_n610), .ZN(
        u4_srl_453_n331) );
  INV_X1 u4_srl_453_U488 ( .A(u4_srl_453_n331), .ZN(u4_srl_453_n596) );
  AOI22_X1 u4_srl_453_U487 ( .A1(u4_srl_453_n20), .A2(u4_srl_453_n505), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n609), .ZN(u4_srl_453_n608) );
  INV_X1 u4_srl_453_U486 ( .A(u4_srl_453_n608), .ZN(u4_srl_453_n607) );
  AOI221_X1 u4_srl_453_U485 ( .B1(u4_srl_453_n506), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n517), .C2(u4_srl_453_n57), .A(u4_srl_453_n607), .ZN(
        u4_srl_453_n310) );
  INV_X1 u4_srl_453_U484 ( .A(u4_srl_453_n310), .ZN(u4_srl_453_n598) );
  INV_X1 u4_srl_453_U483 ( .A(u4_srl_453_n606), .ZN(u4_srl_453_n497) );
  AOI22_X1 u4_srl_453_U482 ( .A1(u4_srl_453_n20), .A2(u4_srl_453_n500), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n605), .ZN(u4_srl_453_n604) );
  OAI221_X1 u4_srl_453_U481 ( .B1(u4_srl_453_n497), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n603), .C2(u4_srl_453_n59), .A(u4_srl_453_n604), .ZN(
        u4_srl_453_n314) );
  INV_X1 u4_srl_453_U480 ( .A(u4_srl_453_n314), .ZN(u4_srl_453_n335) );
  OAI22_X1 u4_srl_453_U479 ( .A1(u4_srl_453_n334), .A2(u4_srl_453_n242), .B1(
        u4_srl_453_n335), .B2(u4_srl_453_n238), .ZN(u4_srl_453_n209) );
  INV_X1 u4_srl_453_U478 ( .A(u4_srl_453_n602), .ZN(u4_srl_453_n492) );
  AOI22_X1 u4_srl_453_U477 ( .A1(u4_srl_453_n20), .A2(u4_srl_453_n495), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n601), .ZN(u4_srl_453_n600) );
  OAI221_X1 u4_srl_453_U476 ( .B1(u4_srl_453_n492), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n599), .C2(u4_srl_453_n59), .A(u4_srl_453_n600), .ZN(
        u4_srl_453_n337) );
  AOI222_X1 u4_srl_453_U475 ( .A1(u4_srl_453_n13), .A2(u4_srl_453_n598), .B1(
        u4_srl_453_n376), .B2(u4_srl_453_n209), .C1(u4_srl_453_n312), .C2(
        u4_srl_453_n337), .ZN(u4_srl_453_n597) );
  OAI221_X1 u4_srl_453_U474 ( .B1(u4_srl_453_n333), .B2(u4_srl_453_n10), .C1(
        u4_srl_453_n596), .C2(u4_srl_453_n8), .A(u4_srl_453_n597), .ZN(
        u4_N5926) );
  AOI22_X1 u4_srl_453_U473 ( .A1(u4_srl_453_n20), .A2(u4_srl_453_n488), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n483), .ZN(u4_srl_453_n595) );
  INV_X1 u4_srl_453_U472 ( .A(u4_srl_453_n595), .ZN(u4_srl_453_n594) );
  AOI221_X1 u4_srl_453_U471 ( .B1(u4_srl_453_n484), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n480), .C2(u4_srl_453_n57), .A(u4_srl_453_n594), .ZN(
        u4_srl_453_n290) );
  AOI22_X1 u4_srl_453_U470 ( .A1(u4_srl_453_n20), .A2(u4_srl_453_n481), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n482), .ZN(u4_srl_453_n593) );
  OAI221_X1 u4_srl_453_U469 ( .B1(u4_srl_453_n478), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n169), .C2(u4_srl_453_n59), .A(u4_srl_453_n593), .ZN(
        u4_srl_453_n287) );
  INV_X1 u4_srl_453_U468 ( .A(u4_srl_453_n287), .ZN(u4_srl_453_n581) );
  AOI22_X1 u4_srl_453_U467 ( .A1(u4_srl_453_n20), .A2(u4_srl_453_n476), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n471), .ZN(u4_srl_453_n592) );
  INV_X1 u4_srl_453_U466 ( .A(u4_srl_453_n592), .ZN(u4_srl_453_n591) );
  AOI221_X1 u4_srl_453_U465 ( .B1(u4_srl_453_n472), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n487), .C2(u4_srl_453_n57), .A(u4_srl_453_n591), .ZN(
        u4_srl_453_n289) );
  INV_X1 u4_srl_453_U464 ( .A(u4_srl_453_n289), .ZN(u4_srl_453_n583) );
  AND2_X1 u4_srl_453_U463 ( .A1(u4_srl_453_n376), .A2(u4_srl_453_n266), .ZN(
        u4_srl_453_n458) );
  AOI22_X1 u4_srl_453_U462 ( .A1(u4_srl_453_n20), .A2(u4_srl_453_n470), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n465), .ZN(u4_srl_453_n590) );
  INV_X1 u4_srl_453_U461 ( .A(u4_srl_453_n590), .ZN(u4_srl_453_n589) );
  AOI221_X1 u4_srl_453_U460 ( .B1(u4_srl_453_n466), .B2(u4_srl_453_n16), .C1(
        u4_srl_453_n462), .C2(u4_srl_453_n57), .A(u4_srl_453_n589), .ZN(
        u4_srl_453_n294) );
  MUX2_X1 u4_srl_453_U459 ( .A(u4_srl_453_n292), .B(u4_srl_453_n294), .S(
        u4_srl_453_n392), .Z(u4_srl_453_n208) );
  INV_X1 u4_srl_453_U458 ( .A(u4_srl_453_n208), .ZN(u4_srl_453_n584) );
  INV_X1 u4_srl_453_U457 ( .A(u4_srl_453_n588), .ZN(u4_srl_453_n460) );
  INV_X1 u4_srl_453_U456 ( .A(u4_srl_453_n475), .ZN(u4_srl_453_n585) );
  AOI22_X1 u4_srl_453_U455 ( .A1(u4_srl_453_n20), .A2(u4_srl_453_n463), .B1(
        u4_srl_453_n28), .B2(u4_srl_453_n587), .ZN(u4_srl_453_n586) );
  OAI221_X1 u4_srl_453_U454 ( .B1(u4_srl_453_n460), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n585), .C2(u4_srl_453_n59), .A(u4_srl_453_n586), .ZN(
        u4_srl_453_n308) );
  AOI222_X1 u4_srl_453_U453 ( .A1(u4_srl_453_n13), .A2(u4_srl_453_n583), .B1(
        u4_srl_453_n458), .B2(u4_srl_453_n584), .C1(u4_srl_453_n312), .C2(
        u4_srl_453_n308), .ZN(u4_srl_453_n582) );
  OAI221_X1 u4_srl_453_U452 ( .B1(u4_srl_453_n290), .B2(u4_srl_453_n9), .C1(
        u4_srl_453_n581), .C2(u4_srl_453_n8), .A(u4_srl_453_n582), .ZN(
        u4_N5927) );
  AOI22_X1 u4_srl_453_U451 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n579), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n580), .ZN(u4_srl_453_n578) );
  INV_X1 u4_srl_453_U450 ( .A(u4_srl_453_n578), .ZN(u4_srl_453_n577) );
  AOI221_X1 u4_srl_453_U449 ( .B1(u4_srl_453_n575), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n576), .C2(u4_srl_453_n57), .A(u4_srl_453_n577), .ZN(
        u4_srl_453_n261) );
  AOI22_X1 u4_srl_453_U448 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n573), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n574), .ZN(u4_srl_453_n572) );
  OAI221_X1 u4_srl_453_U447 ( .B1(u4_srl_453_n570), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n571), .C2(u4_srl_453_n58), .A(u4_srl_453_n572), .ZN(
        u4_srl_453_n258) );
  INV_X1 u4_srl_453_U446 ( .A(u4_srl_453_n258), .ZN(u4_srl_453_n550) );
  AOI22_X1 u4_srl_453_U445 ( .A1(u4_srl_453_n20), .A2(u4_srl_453_n568), .B1(
        u4_srl_453_n25), .B2(u4_srl_453_n569), .ZN(u4_srl_453_n567) );
  INV_X1 u4_srl_453_U444 ( .A(u4_srl_453_n567), .ZN(u4_srl_453_n566) );
  AOI221_X1 u4_srl_453_U443 ( .B1(u4_srl_453_n564), .B2(u4_srl_453_n15), .C1(
        u4_srl_453_n565), .C2(u4_srl_453_n57), .A(u4_srl_453_n566), .ZN(
        u4_srl_453_n260) );
  INV_X1 u4_srl_453_U442 ( .A(u4_srl_453_n260), .ZN(u4_srl_453_n552) );
  AOI22_X1 u4_srl_453_U441 ( .A1(u4_srl_453_n394), .A2(u4_srl_453_n562), .B1(
        u4_srl_453_n25), .B2(u4_srl_453_n563), .ZN(u4_srl_453_n561) );
  INV_X1 u4_srl_453_U440 ( .A(u4_srl_453_n561), .ZN(u4_srl_453_n560) );
  AOI221_X1 u4_srl_453_U439 ( .B1(u4_srl_453_n558), .B2(u4_srl_453_n15), .C1(
        u4_srl_453_n559), .C2(u4_srl_453_n409), .A(u4_srl_453_n560), .ZN(
        u4_srl_453_n264) );
  NAND2_X1 u4_srl_453_U438 ( .A1(u4_srl_453_n409), .A2(u4_shift_right[4]), 
        .ZN(u4_srl_453_n464) );
  OAI22_X1 u4_srl_453_U437 ( .A1(u4_shift_right[4]), .A2(u4_srl_453_n264), 
        .B1(u4_srl_453_n263), .B2(u4_srl_453_n464), .ZN(u4_srl_453_n306) );
  AOI22_X1 u4_srl_453_U436 ( .A1(u4_srl_453_n20), .A2(u4_srl_453_n556), .B1(
        u4_srl_453_n28), .B2(u4_srl_453_n557), .ZN(u4_srl_453_n555) );
  OAI221_X1 u4_srl_453_U435 ( .B1(u4_srl_453_n553), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n554), .C2(u4_srl_453_n59), .A(u4_srl_453_n555), .ZN(
        u4_srl_453_n307) );
  AOI222_X1 u4_srl_453_U434 ( .A1(u4_srl_453_n13), .A2(u4_srl_453_n552), .B1(
        u4_srl_453_n458), .B2(u4_srl_453_n306), .C1(u4_srl_453_n312), .C2(
        u4_srl_453_n307), .ZN(u4_srl_453_n551) );
  OAI221_X1 u4_srl_453_U433 ( .B1(u4_srl_453_n261), .B2(u4_srl_453_n10), .C1(
        u4_srl_453_n550), .C2(u4_srl_453_n8), .A(u4_srl_453_n551), .ZN(
        u4_N5928) );
  AOI22_X1 u4_srl_453_U432 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n548), .B1(
        u4_srl_453_n28), .B2(u4_srl_453_n549), .ZN(u4_srl_453_n547) );
  INV_X1 u4_srl_453_U431 ( .A(u4_srl_453_n547), .ZN(u4_srl_453_n546) );
  AOI221_X1 u4_srl_453_U430 ( .B1(u4_srl_453_n544), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n545), .C2(u4_srl_453_n57), .A(u4_srl_453_n546), .ZN(
        u4_srl_453_n230) );
  AOI22_X1 u4_srl_453_U429 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n542), .B1(
        u4_srl_453_n28), .B2(u4_srl_453_n543), .ZN(u4_srl_453_n541) );
  OAI221_X1 u4_srl_453_U428 ( .B1(u4_srl_453_n539), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n540), .C2(u4_srl_453_n59), .A(u4_srl_453_n541), .ZN(
        u4_srl_453_n226) );
  INV_X1 u4_srl_453_U427 ( .A(u4_srl_453_n226), .ZN(u4_srl_453_n519) );
  AOI22_X1 u4_srl_453_U426 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n537), .B1(
        u4_srl_453_n25), .B2(u4_srl_453_n538), .ZN(u4_srl_453_n536) );
  INV_X1 u4_srl_453_U425 ( .A(u4_srl_453_n536), .ZN(u4_srl_453_n535) );
  AOI221_X1 u4_srl_453_U424 ( .B1(u4_srl_453_n533), .B2(u4_srl_453_n15), .C1(
        u4_srl_453_n534), .C2(u4_srl_453_n56), .A(u4_srl_453_n535), .ZN(
        u4_srl_453_n229) );
  INV_X1 u4_srl_453_U423 ( .A(u4_srl_453_n229), .ZN(u4_srl_453_n521) );
  AOI22_X1 u4_srl_453_U422 ( .A1(u4_srl_453_n394), .A2(u4_srl_453_n531), .B1(
        u4_srl_453_n25), .B2(u4_srl_453_n532), .ZN(u4_srl_453_n530) );
  INV_X1 u4_srl_453_U421 ( .A(u4_srl_453_n530), .ZN(u4_srl_453_n529) );
  AOI221_X1 u4_srl_453_U420 ( .B1(u4_srl_453_n527), .B2(u4_srl_453_n15), .C1(
        u4_srl_453_n528), .C2(u4_srl_453_n56), .A(u4_srl_453_n529), .ZN(
        u4_srl_453_n248) );
  OAI22_X1 u4_srl_453_U419 ( .A1(u4_shift_right[4]), .A2(u4_srl_453_n248), 
        .B1(u4_srl_453_n247), .B2(u4_srl_453_n464), .ZN(u4_srl_453_n304) );
  AOI22_X1 u4_srl_453_U418 ( .A1(u4_srl_453_n22), .A2(u4_srl_453_n525), .B1(
        u4_srl_453_n28), .B2(u4_srl_453_n526), .ZN(u4_srl_453_n524) );
  OAI221_X1 u4_srl_453_U417 ( .B1(u4_srl_453_n522), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n523), .C2(u4_srl_453_n59), .A(u4_srl_453_n524), .ZN(
        u4_srl_453_n305) );
  AOI222_X1 u4_srl_453_U416 ( .A1(u4_srl_453_n13), .A2(u4_srl_453_n521), .B1(
        u4_srl_453_n458), .B2(u4_srl_453_n304), .C1(u4_srl_453_n312), .C2(
        u4_srl_453_n305), .ZN(u4_srl_453_n520) );
  OAI221_X1 u4_srl_453_U415 ( .B1(u4_srl_453_n230), .B2(u4_srl_453_n9), .C1(
        u4_srl_453_n519), .C2(u4_srl_453_n8), .A(u4_srl_453_n520), .ZN(
        u4_N5929) );
  AOI22_X1 u4_srl_453_U414 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n517), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n518), .ZN(u4_srl_453_n516) );
  INV_X1 u4_srl_453_U413 ( .A(u4_srl_453_n516), .ZN(u4_srl_453_n515) );
  AOI221_X1 u4_srl_453_U412 ( .B1(u4_srl_453_n513), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n514), .C2(u4_srl_453_n56), .A(u4_srl_453_n515), .ZN(
        u4_srl_453_n202) );
  INV_X1 u4_srl_453_U411 ( .A(u4_srl_453_n512), .ZN(u4_srl_453_n507) );
  AOI22_X1 u4_srl_453_U410 ( .A1(u4_srl_453_n22), .A2(u4_srl_453_n510), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n511), .ZN(u4_srl_453_n509) );
  OAI221_X1 u4_srl_453_U409 ( .B1(u4_srl_453_n507), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n508), .C2(u4_srl_453_n59), .A(u4_srl_453_n509), .ZN(
        u4_srl_453_n198) );
  INV_X1 u4_srl_453_U408 ( .A(u4_srl_453_n198), .ZN(u4_srl_453_n489) );
  INV_X1 u4_srl_453_U407 ( .A(u4_srl_453_n506), .ZN(u4_srl_453_n502) );
  AOI22_X1 u4_srl_453_U406 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n504), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n505), .ZN(u4_srl_453_n503) );
  OAI221_X1 u4_srl_453_U405 ( .B1(u4_srl_453_n501), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n502), .C2(u4_srl_453_n59), .A(u4_srl_453_n503), .ZN(
        u4_srl_453_n382) );
  AOI22_X1 u4_srl_453_U404 ( .A1(u4_srl_453_n23), .A2(u4_srl_453_n499), .B1(
        u4_srl_453_n27), .B2(u4_srl_453_n500), .ZN(u4_srl_453_n498) );
  OAI221_X1 u4_srl_453_U403 ( .B1(u4_srl_453_n496), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n497), .C2(u4_srl_453_n59), .A(u4_srl_453_n498), .ZN(
        u4_srl_453_n381) );
  INV_X1 u4_srl_453_U402 ( .A(u4_srl_453_n381), .ZN(u4_srl_453_n245) );
  OAI22_X1 u4_srl_453_U401 ( .A1(u4_shift_right[4]), .A2(u4_srl_453_n245), 
        .B1(u4_srl_453_n244), .B2(u4_srl_453_n464), .ZN(u4_srl_453_n302) );
  AOI22_X1 u4_srl_453_U400 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n494), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n495), .ZN(u4_srl_453_n493) );
  OAI221_X1 u4_srl_453_U399 ( .B1(u4_srl_453_n491), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n492), .C2(u4_srl_453_n59), .A(u4_srl_453_n493), .ZN(
        u4_srl_453_n303) );
  AOI222_X1 u4_srl_453_U398 ( .A1(u4_srl_453_n13), .A2(u4_srl_453_n382), .B1(
        u4_srl_453_n458), .B2(u4_srl_453_n302), .C1(u4_srl_453_n312), .C2(
        u4_srl_453_n303), .ZN(u4_srl_453_n490) );
  OAI221_X1 u4_srl_453_U397 ( .B1(u4_srl_453_n202), .B2(u4_srl_453_n10), .C1(
        u4_srl_453_n489), .C2(u4_srl_453_n8), .A(u4_srl_453_n490), .ZN(
        u4_N5930) );
  AOI22_X1 u4_srl_453_U396 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n487), .B1(
        u4_srl_453_n26), .B2(u4_srl_453_n488), .ZN(u4_srl_453_n486) );
  INV_X1 u4_srl_453_U395 ( .A(u4_srl_453_n486), .ZN(u4_srl_453_n485) );
  AOI221_X1 u4_srl_453_U394 ( .B1(u4_srl_453_n483), .B2(u4_srl_453_n15), .C1(
        u4_srl_453_n484), .C2(u4_srl_453_n56), .A(u4_srl_453_n485), .ZN(
        u4_srl_453_n178) );
  INV_X1 u4_srl_453_U393 ( .A(u4_srl_453_n482), .ZN(u4_srl_453_n477) );
  AOI22_X1 u4_srl_453_U392 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n480), .B1(
        u4_srl_453_n25), .B2(u4_srl_453_n481), .ZN(u4_srl_453_n479) );
  OAI221_X1 u4_srl_453_U391 ( .B1(u4_srl_453_n477), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n478), .C2(u4_srl_453_n59), .A(u4_srl_453_n479), .ZN(
        u4_srl_453_n172) );
  INV_X1 u4_srl_453_U390 ( .A(u4_srl_453_n172), .ZN(u4_srl_453_n455) );
  AOI22_X1 u4_srl_453_U389 ( .A1(u4_srl_453_n21), .A2(u4_srl_453_n475), .B1(
        u4_srl_453_n25), .B2(u4_srl_453_n476), .ZN(u4_srl_453_n474) );
  INV_X1 u4_srl_453_U388 ( .A(u4_srl_453_n474), .ZN(u4_srl_453_n473) );
  AOI221_X1 u4_srl_453_U387 ( .B1(u4_srl_453_n471), .B2(u4_srl_453_n17), .C1(
        u4_srl_453_n472), .C2(u4_srl_453_n56), .A(u4_srl_453_n473), .ZN(
        u4_srl_453_n176) );
  INV_X1 u4_srl_453_U386 ( .A(u4_srl_453_n176), .ZN(u4_srl_453_n457) );
  AOI22_X1 u4_srl_453_U385 ( .A1(u4_srl_453_n22), .A2(u4_srl_453_n469), .B1(
        u4_srl_453_n28), .B2(u4_srl_453_n470), .ZN(u4_srl_453_n468) );
  INV_X1 u4_srl_453_U384 ( .A(u4_srl_453_n468), .ZN(u4_srl_453_n467) );
  AOI221_X1 u4_srl_453_U383 ( .B1(u4_srl_453_n465), .B2(u4_srl_453_n15), .C1(
        u4_srl_453_n466), .C2(u4_srl_453_n56), .A(u4_srl_453_n467), .ZN(
        u4_srl_453_n241) );
  OAI22_X1 u4_srl_453_U382 ( .A1(u4_srl_453_n241), .A2(u4_shift_right[4]), 
        .B1(u4_srl_453_n240), .B2(u4_srl_453_n464), .ZN(u4_srl_453_n300) );
  AOI22_X1 u4_srl_453_U381 ( .A1(u4_srl_453_n20), .A2(u4_srl_453_n462), .B1(
        u4_srl_453_n25), .B2(u4_srl_453_n463), .ZN(u4_srl_453_n461) );
  OAI221_X1 u4_srl_453_U380 ( .B1(u4_srl_453_n459), .B2(u4_srl_453_n18), .C1(
        u4_srl_453_n460), .C2(u4_srl_453_n59), .A(u4_srl_453_n461), .ZN(
        u4_srl_453_n301) );
  AOI222_X1 u4_srl_453_U379 ( .A1(u4_srl_453_n13), .A2(u4_srl_453_n457), .B1(
        u4_srl_453_n458), .B2(u4_srl_453_n300), .C1(u4_srl_453_n312), .C2(
        u4_srl_453_n301), .ZN(u4_srl_453_n456) );
  OAI221_X1 u4_srl_453_U378 ( .B1(u4_srl_453_n178), .B2(u4_srl_453_n10), .C1(
        u4_srl_453_n455), .C2(u4_srl_453_n8), .A(u4_srl_453_n456), .ZN(
        u4_N5931) );
  INV_X1 u4_srl_453_U377 ( .A(u4_srl_453_n298), .ZN(u4_srl_453_n454) );
  INV_X1 u4_srl_453_U376 ( .A(u4_srl_453_n190), .ZN(u4_srl_453_n370) );
  AOI222_X1 u4_srl_453_U375 ( .A1(u4_srl_453_n13), .A2(u4_srl_453_n454), .B1(
        u4_srl_453_n12), .B2(u4_srl_453_n371), .C1(u4_srl_453_n408), .C2(
        u4_srl_453_n370), .ZN(u4_srl_453_n453) );
  OAI221_X1 u4_srl_453_U374 ( .B1(u4_srl_453_n373), .B2(u4_srl_453_n10), .C1(
        u4_srl_453_n452), .C2(u4_srl_453_n8), .A(u4_srl_453_n453), .ZN(
        u4_N5932) );
  INV_X1 u4_srl_453_U373 ( .A(u4_srl_453_n296), .ZN(u4_srl_453_n451) );
  INV_X1 u4_srl_453_U372 ( .A(u4_srl_453_n189), .ZN(u4_srl_453_n365) );
  AOI222_X1 u4_srl_453_U371 ( .A1(u4_srl_453_n13), .A2(u4_srl_453_n451), .B1(
        u4_srl_453_n12), .B2(u4_srl_453_n366), .C1(u4_srl_453_n408), .C2(
        u4_srl_453_n365), .ZN(u4_srl_453_n450) );
  OAI221_X1 u4_srl_453_U370 ( .B1(u4_srl_453_n368), .B2(u4_srl_453_n10), .C1(
        u4_srl_453_n449), .C2(u4_srl_453_n8), .A(u4_srl_453_n450), .ZN(
        u4_N5933) );
  AOI222_X1 u4_srl_453_U369 ( .A1(u4_srl_453_n13), .A2(u4_srl_453_n448), .B1(
        u4_srl_453_n12), .B2(u4_srl_453_n361), .C1(u4_srl_453_n408), .C2(
        u4_srl_453_n360), .ZN(u4_srl_453_n447) );
  OAI221_X1 u4_srl_453_U368 ( .B1(u4_srl_453_n363), .B2(u4_srl_453_n10), .C1(
        u4_srl_453_n446), .C2(u4_srl_453_n8), .A(u4_srl_453_n447), .ZN(
        u4_N5934) );
  INV_X1 u4_srl_453_U367 ( .A(u4_srl_453_n278), .ZN(u4_srl_453_n445) );
  INV_X1 u4_srl_453_U366 ( .A(u4_srl_453_n187), .ZN(u4_srl_453_n355) );
  AOI222_X1 u4_srl_453_U365 ( .A1(u4_srl_453_n13), .A2(u4_srl_453_n445), .B1(
        u4_srl_453_n12), .B2(u4_srl_453_n356), .C1(u4_srl_453_n408), .C2(
        u4_srl_453_n355), .ZN(u4_srl_453_n444) );
  OAI221_X1 u4_srl_453_U364 ( .B1(u4_srl_453_n358), .B2(u4_srl_453_n10), .C1(
        u4_srl_453_n443), .C2(u4_srl_453_n8), .A(u4_srl_453_n444), .ZN(
        u4_N5935) );
  AOI222_X1 u4_srl_453_U363 ( .A1(u4_srl_453_n417), .A2(u4_srl_453_n400), .B1(
        u4_srl_453_n323), .B2(u4_srl_453_n336), .C1(u4_srl_453_n324), .C2(
        u4_srl_453_n401), .ZN(u4_srl_453_n270) );
  INV_X1 u4_srl_453_U362 ( .A(u4_srl_453_n415), .ZN(u4_srl_453_n435) );
  OAI22_X1 u4_srl_453_U361 ( .A1(u4_srl_453_n36), .A2(u4_srl_453_n60), .B1(
        u4_srl_453_n29), .B2(u4_srl_453_n61), .ZN(u4_srl_453_n442) );
  AOI221_X1 u4_srl_453_U360 ( .B1(n6348), .B2(u4_srl_453_n42), .C1(n6347), 
        .C2(u4_srl_453_n47), .A(u4_srl_453_n442), .ZN(u4_srl_453_n437) );
  AOI22_X1 u4_srl_453_U359 ( .A1(n6444), .A2(u4_srl_453_n42), .B1(n6351), .B2(
        u4_srl_453_n47), .ZN(u4_srl_453_n441) );
  OAI221_X1 u4_srl_453_U358 ( .B1(u4_srl_453_n29), .B2(u4_srl_453_n65), .C1(
        u4_srl_453_n36), .C2(u4_srl_453_n64), .A(u4_srl_453_n441), .ZN(
        u4_srl_453_n256) );
  AOI222_X1 u4_srl_453_U357 ( .A1(u4_srl_453_n15), .A2(u4_srl_453_n256), .B1(
        u4_srl_453_n21), .B2(u4_srl_453_n253), .C1(u4_srl_453_n25), .C2(
        u4_srl_453_n257), .ZN(u4_srl_453_n440) );
  MUX2_X1 u4_srl_453_U356 ( .A(u4_srl_453_n439), .B(u4_srl_453_n440), .S(
        u4_srl_453_n392), .Z(u4_srl_453_n438) );
  OAI21_X1 u4_srl_453_U355 ( .B1(u4_srl_453_n437), .B2(u4_srl_453_n265), .A(
        u4_srl_453_n438), .ZN(u4_srl_453_n436) );
  AOI22_X1 u4_srl_453_U354 ( .A1(u4_srl_453_n14), .A2(u4_srl_453_n435), .B1(
        u4_srl_453_n386), .B2(u4_srl_453_n436), .ZN(u4_srl_453_n434) );
  OAI221_X1 u4_srl_453_U353 ( .B1(u4_srl_453_n270), .B2(u4_srl_453_n383), .C1(
        u4_srl_453_n321), .C2(u4_srl_453_n11), .A(u4_srl_453_n434), .ZN(
        u4_N5908) );
  INV_X1 u4_srl_453_U352 ( .A(u4_srl_453_n276), .ZN(u4_srl_453_n431) );
  INV_X1 u4_srl_453_U351 ( .A(u4_srl_453_n186), .ZN(u4_srl_453_n433) );
  AOI222_X1 u4_srl_453_U350 ( .A1(u4_srl_453_n13), .A2(u4_srl_453_n431), .B1(
        u4_srl_453_n12), .B2(u4_srl_453_n432), .C1(u4_srl_453_n408), .C2(
        u4_srl_453_n433), .ZN(u4_srl_453_n430) );
  OAI221_X1 u4_srl_453_U349 ( .B1(u4_srl_453_n353), .B2(u4_srl_453_n10), .C1(
        u4_srl_453_n429), .C2(u4_srl_453_n8), .A(u4_srl_453_n430), .ZN(
        u4_N5936) );
  INV_X1 u4_srl_453_U348 ( .A(u4_srl_453_n185), .ZN(u4_srl_453_n428) );
  AOI222_X1 u4_srl_453_U347 ( .A1(u4_srl_453_n14), .A2(u4_srl_453_n426), .B1(
        u4_srl_453_n12), .B2(u4_srl_453_n427), .C1(u4_srl_453_n408), .C2(
        u4_srl_453_n428), .ZN(u4_srl_453_n425) );
  OAI221_X1 u4_srl_453_U346 ( .B1(u4_srl_453_n350), .B2(u4_srl_453_n9), .C1(
        u4_srl_453_n424), .C2(u4_srl_453_n8), .A(u4_srl_453_n425), .ZN(
        u4_N5937) );
  AOI222_X1 u4_srl_453_U345 ( .A1(u4_srl_453_n13), .A2(u4_srl_453_n423), .B1(
        u4_srl_453_n12), .B2(u4_srl_453_n347), .C1(u4_srl_453_n408), .C2(
        u4_srl_453_n346), .ZN(u4_srl_453_n422) );
  OAI221_X1 u4_srl_453_U344 ( .B1(u4_srl_453_n344), .B2(u4_srl_453_n9), .C1(
        u4_srl_453_n421), .C2(u4_srl_453_n8), .A(u4_srl_453_n422), .ZN(
        u4_N5938) );
  AOI222_X1 u4_srl_453_U343 ( .A1(u4_srl_453_n14), .A2(u4_srl_453_n420), .B1(
        u4_srl_453_n12), .B2(u4_srl_453_n342), .C1(u4_srl_453_n408), .C2(
        u4_srl_453_n341), .ZN(u4_srl_453_n419) );
  OAI221_X1 u4_srl_453_U342 ( .B1(u4_srl_453_n339), .B2(u4_srl_453_n9), .C1(
        u4_srl_453_n418), .C2(u4_srl_453_n8), .A(u4_srl_453_n419), .ZN(
        u4_N5939) );
  AOI222_X1 u4_srl_453_U341 ( .A1(u4_srl_453_n14), .A2(u4_srl_453_n417), .B1(
        u4_srl_453_n12), .B2(u4_srl_453_n324), .C1(u4_srl_453_n408), .C2(
        u4_srl_453_n323), .ZN(u4_srl_453_n416) );
  OAI221_X1 u4_srl_453_U340 ( .B1(u4_srl_453_n321), .B2(u4_srl_453_n9), .C1(
        u4_srl_453_n415), .C2(u4_srl_453_n8), .A(u4_srl_453_n416), .ZN(
        u4_N5940) );
  AOI222_X1 u4_srl_453_U339 ( .A1(u4_srl_453_n13), .A2(u4_srl_453_n399), .B1(
        u4_srl_453_n12), .B2(u4_srl_453_n319), .C1(u4_srl_453_n408), .C2(
        u4_srl_453_n318), .ZN(u4_srl_453_n414) );
  OAI221_X1 u4_srl_453_U338 ( .B1(u4_srl_453_n316), .B2(u4_srl_453_n9), .C1(
        u4_srl_453_n398), .C2(u4_srl_453_n8), .A(u4_srl_453_n414), .ZN(
        u4_N5941) );
  INV_X1 u4_srl_453_U337 ( .A(u4_srl_453_n334), .ZN(u4_srl_453_n313) );
  AOI222_X1 u4_srl_453_U336 ( .A1(u4_srl_453_n13), .A2(u4_srl_453_n337), .B1(
        u4_srl_453_n12), .B2(u4_srl_453_n314), .C1(u4_srl_453_n408), .C2(
        u4_srl_453_n313), .ZN(u4_srl_453_n413) );
  OAI221_X1 u4_srl_453_U335 ( .B1(u4_srl_453_n310), .B2(u4_srl_453_n9), .C1(
        u4_srl_453_n333), .C2(u4_srl_453_n8), .A(u4_srl_453_n413), .ZN(
        u4_N5942) );
  INV_X1 u4_srl_453_U334 ( .A(u4_srl_453_n292), .ZN(u4_srl_453_n411) );
  INV_X1 u4_srl_453_U333 ( .A(u4_srl_453_n294), .ZN(u4_srl_453_n412) );
  AOI222_X1 u4_srl_453_U332 ( .A1(u4_srl_453_n14), .A2(u4_srl_453_n308), .B1(
        u4_srl_453_n408), .B2(u4_srl_453_n411), .C1(u4_srl_453_n12), .C2(
        u4_srl_453_n412), .ZN(u4_srl_453_n410) );
  OAI221_X1 u4_srl_453_U331 ( .B1(u4_srl_453_n289), .B2(u4_srl_453_n9), .C1(
        u4_srl_453_n290), .C2(u4_srl_453_n8), .A(u4_srl_453_n410), .ZN(
        u4_N5943) );
  AND2_X1 u4_srl_453_U330 ( .A1(u4_srl_453_n408), .A2(u4_srl_453_n409), .ZN(
        u4_srl_453_n379) );
  INV_X1 u4_srl_453_U329 ( .A(u4_srl_453_n264), .ZN(u4_srl_453_n407) );
  AOI222_X1 u4_srl_453_U328 ( .A1(u4_srl_453_n14), .A2(u4_srl_453_n307), .B1(
        u4_srl_453_n379), .B2(u4_srl_453_n406), .C1(u4_srl_453_n12), .C2(
        u4_srl_453_n407), .ZN(u4_srl_453_n405) );
  OAI221_X1 u4_srl_453_U327 ( .B1(u4_srl_453_n260), .B2(u4_srl_453_n9), .C1(
        u4_srl_453_n261), .C2(u4_srl_453_n8), .A(u4_srl_453_n405), .ZN(
        u4_N5944) );
  INV_X1 u4_srl_453_U326 ( .A(u4_srl_453_n248), .ZN(u4_srl_453_n404) );
  AOI222_X1 u4_srl_453_U325 ( .A1(u4_srl_453_n13), .A2(u4_srl_453_n305), .B1(
        u4_srl_453_n379), .B2(u4_srl_453_n403), .C1(u4_srl_453_n12), .C2(
        u4_srl_453_n404), .ZN(u4_srl_453_n402) );
  OAI221_X1 u4_srl_453_U324 ( .B1(u4_srl_453_n229), .B2(u4_srl_453_n9), .C1(
        u4_srl_453_n230), .C2(u4_srl_453_n8), .A(u4_srl_453_n402), .ZN(
        u4_N5945) );
  AOI222_X1 u4_srl_453_U323 ( .A1(u4_srl_453_n399), .A2(u4_srl_453_n400), .B1(
        u4_srl_453_n318), .B2(u4_srl_453_n336), .C1(u4_srl_453_n319), .C2(
        u4_srl_453_n401), .ZN(u4_srl_453_n269) );
  INV_X1 u4_srl_453_U322 ( .A(u4_srl_453_n398), .ZN(u4_srl_453_n385) );
  OAI22_X1 u4_srl_453_U321 ( .A1(u4_srl_453_n36), .A2(u4_srl_453_n61), .B1(
        u4_srl_453_n29), .B2(u4_srl_453_n62), .ZN(u4_srl_453_n397) );
  AOI221_X1 u4_srl_453_U320 ( .B1(n6349), .B2(u4_srl_453_n42), .C1(n6348), 
        .C2(u4_srl_453_n47), .A(u4_srl_453_n397), .ZN(u4_srl_453_n388) );
  AOI22_X1 u4_srl_453_U319 ( .A1(n6443), .A2(u4_srl_453_n44), .B1(n6444), .B2(
        u4_srl_453_n47), .ZN(u4_srl_453_n395) );
  OAI221_X1 u4_srl_453_U318 ( .B1(u4_srl_453_n31), .B2(u4_srl_453_n66), .C1(
        u4_srl_453_n39), .C2(u4_srl_453_n65), .A(u4_srl_453_n395), .ZN(
        u4_srl_453_n224) );
  AOI222_X1 u4_srl_453_U317 ( .A1(u4_srl_453_n15), .A2(u4_srl_453_n224), .B1(
        u4_srl_453_n21), .B2(u4_srl_453_n221), .C1(u4_srl_453_n25), .C2(
        u4_srl_453_n225), .ZN(u4_srl_453_n391) );
  MUX2_X1 u4_srl_453_U316 ( .A(u4_srl_453_n390), .B(u4_srl_453_n391), .S(
        u4_srl_453_n392), .Z(u4_srl_453_n389) );
  OAI21_X1 u4_srl_453_U315 ( .B1(u4_srl_453_n388), .B2(u4_srl_453_n265), .A(
        u4_srl_453_n389), .ZN(u4_srl_453_n387) );
  AOI22_X1 u4_srl_453_U314 ( .A1(u4_srl_453_n14), .A2(u4_srl_453_n385), .B1(
        u4_srl_453_n386), .B2(u4_srl_453_n387), .ZN(u4_srl_453_n384) );
  OAI221_X1 u4_srl_453_U313 ( .B1(u4_srl_453_n269), .B2(u4_srl_453_n383), .C1(
        u4_srl_453_n316), .C2(u4_srl_453_n11), .A(u4_srl_453_n384), .ZN(
        u4_N5909) );
  INV_X1 u4_srl_453_U312 ( .A(u4_srl_453_n382), .ZN(u4_srl_453_n201) );
  AOI222_X1 u4_srl_453_U311 ( .A1(u4_srl_453_n13), .A2(u4_srl_453_n303), .B1(
        u4_srl_453_n379), .B2(u4_srl_453_n380), .C1(u4_srl_453_n12), .C2(
        u4_srl_453_n381), .ZN(u4_srl_453_n378) );
  OAI221_X1 u4_srl_453_U310 ( .B1(u4_srl_453_n201), .B2(u4_srl_453_n9), .C1(
        u4_srl_453_n202), .C2(u4_srl_453_n8), .A(u4_srl_453_n378), .ZN(
        u4_N5946) );
  INV_X1 u4_srl_453_U309 ( .A(u4_srl_453_n241), .ZN(u4_srl_453_n377) );
  AOI222_X1 u4_srl_453_U308 ( .A1(u4_srl_453_n14), .A2(u4_srl_453_n301), .B1(
        u4_srl_453_n375), .B2(u4_srl_453_n376), .C1(u4_srl_453_n312), .C2(
        u4_srl_453_n377), .ZN(u4_srl_453_n374) );
  OAI221_X1 u4_srl_453_U307 ( .B1(u4_srl_453_n176), .B2(u4_srl_453_n9), .C1(
        u4_srl_453_n178), .C2(u4_srl_453_n8), .A(u4_srl_453_n374), .ZN(
        u4_N5947) );
  OAI22_X1 u4_srl_453_U306 ( .A1(u4_srl_453_n9), .A2(u4_srl_453_n298), .B1(
        u4_srl_453_n8), .B2(u4_srl_453_n373), .ZN(u4_srl_453_n372) );
  AOI221_X1 u4_srl_453_U305 ( .B1(u4_srl_453_n370), .B2(u4_srl_453_n312), .C1(
        u4_srl_453_n371), .C2(u4_srl_453_n14), .A(u4_srl_453_n372), .ZN(
        u4_srl_453_n369) );
  INV_X1 u4_srl_453_U304 ( .A(u4_srl_453_n369), .ZN(u4_N5948) );
  OAI22_X1 u4_srl_453_U303 ( .A1(u4_srl_453_n10), .A2(u4_srl_453_n296), .B1(
        u4_srl_453_n8), .B2(u4_srl_453_n368), .ZN(u4_srl_453_n367) );
  AOI221_X1 u4_srl_453_U302 ( .B1(u4_srl_453_n365), .B2(u4_srl_453_n312), .C1(
        u4_srl_453_n366), .C2(u4_srl_453_n14), .A(u4_srl_453_n367), .ZN(
        u4_srl_453_n364) );
  INV_X1 u4_srl_453_U301 ( .A(u4_srl_453_n364), .ZN(u4_N5949) );
  OAI22_X1 u4_srl_453_U300 ( .A1(u4_srl_453_n9), .A2(u4_srl_453_n280), .B1(
        u4_srl_453_n8), .B2(u4_srl_453_n363), .ZN(u4_srl_453_n362) );
  AOI221_X1 u4_srl_453_U299 ( .B1(u4_srl_453_n360), .B2(u4_srl_453_n312), .C1(
        u4_srl_453_n361), .C2(u4_srl_453_n14), .A(u4_srl_453_n362), .ZN(
        u4_srl_453_n359) );
  INV_X1 u4_srl_453_U298 ( .A(u4_srl_453_n359), .ZN(u4_N5950) );
  OAI22_X1 u4_srl_453_U297 ( .A1(u4_srl_453_n9), .A2(u4_srl_453_n278), .B1(
        u4_srl_453_n8), .B2(u4_srl_453_n358), .ZN(u4_srl_453_n357) );
  AOI221_X1 u4_srl_453_U296 ( .B1(u4_srl_453_n355), .B2(u4_srl_453_n312), .C1(
        u4_srl_453_n356), .C2(u4_srl_453_n14), .A(u4_srl_453_n357), .ZN(
        u4_srl_453_n354) );
  INV_X1 u4_srl_453_U295 ( .A(u4_srl_453_n354), .ZN(u4_N5951) );
  OAI22_X1 u4_srl_453_U294 ( .A1(u4_srl_453_n9), .A2(u4_srl_453_n276), .B1(
        u4_srl_453_n8), .B2(u4_srl_453_n353), .ZN(u4_srl_453_n352) );
  INV_X1 u4_srl_453_U293 ( .A(u4_srl_453_n352), .ZN(u4_srl_453_n351) );
  OAI221_X1 u4_srl_453_U292 ( .B1(u4_srl_453_n186), .B2(u4_srl_453_n11), .C1(
        u4_srl_453_n275), .C2(u4_srl_453_n4), .A(u4_srl_453_n351), .ZN(
        u4_N5952) );
  OAI22_X1 u4_srl_453_U291 ( .A1(u4_srl_453_n9), .A2(u4_srl_453_n274), .B1(
        u4_srl_453_n8), .B2(u4_srl_453_n350), .ZN(u4_srl_453_n349) );
  INV_X1 u4_srl_453_U290 ( .A(u4_srl_453_n349), .ZN(u4_srl_453_n348) );
  OAI221_X1 u4_srl_453_U289 ( .B1(u4_srl_453_n185), .B2(u4_srl_453_n11), .C1(
        u4_srl_453_n273), .C2(u4_srl_453_n4), .A(u4_srl_453_n348), .ZN(
        u4_N5953) );
  AOI22_X1 u4_srl_453_U288 ( .A1(u4_srl_453_n12), .A2(u4_srl_453_n346), .B1(
        u4_srl_453_n14), .B2(u4_srl_453_n347), .ZN(u4_srl_453_n345) );
  OAI221_X1 u4_srl_453_U287 ( .B1(u4_srl_453_n343), .B2(u4_srl_453_n9), .C1(
        u4_srl_453_n344), .C2(u4_srl_453_n8), .A(u4_srl_453_n345), .ZN(
        u4_N5954) );
  AOI22_X1 u4_srl_453_U286 ( .A1(u4_srl_453_n12), .A2(u4_srl_453_n341), .B1(
        u4_srl_453_n14), .B2(u4_srl_453_n342), .ZN(u4_srl_453_n340) );
  OAI221_X1 u4_srl_453_U285 ( .B1(u4_srl_453_n338), .B2(u4_srl_453_n9), .C1(
        u4_srl_453_n339), .C2(u4_srl_453_n8), .A(u4_srl_453_n340), .ZN(
        u4_N5955) );
  INV_X1 u4_srl_453_U284 ( .A(u4_srl_453_n337), .ZN(u4_srl_453_n309) );
  INV_X1 u4_srl_453_U283 ( .A(u4_srl_453_n336), .ZN(u4_srl_453_n293) );
  OAI222_X1 u4_srl_453_U282 ( .A1(u4_srl_453_n309), .A2(u4_srl_453_n238), .B1(
        u4_srl_453_n334), .B2(u4_srl_453_n293), .C1(u4_srl_453_n335), .C2(
        u4_srl_453_n242), .ZN(u4_srl_453_n268) );
  OAI22_X1 u4_srl_453_U281 ( .A1(u4_srl_453_n310), .A2(u4_srl_453_n177), .B1(
        u4_srl_453_n333), .B2(u4_srl_453_n179), .ZN(u4_srl_453_n332) );
  AOI221_X1 u4_srl_453_U280 ( .B1(u4_srl_453_n171), .B2(u4_srl_453_n331), .C1(
        u4_srl_453_n268), .C2(u4_srl_453_n174), .A(u4_srl_453_n332), .ZN(
        u4_srl_453_n325) );
  INV_X1 u4_srl_453_U279 ( .A(u4_srl_453_n170), .ZN(u4_srl_453_n218) );
  INV_X1 u4_srl_453_U278 ( .A(u4_srl_453_n168), .ZN(u4_srl_453_n220) );
  AOI22_X1 u4_srl_453_U277 ( .A1(u4_srl_453_n330), .A2(u4_srl_453_n164), .B1(
        u4_srl_453_n194), .B2(u4_srl_453_n162), .ZN(u4_srl_453_n329) );
  INV_X1 u4_srl_453_U276 ( .A(u4_srl_453_n329), .ZN(u4_srl_453_n328) );
  AOI221_X1 u4_srl_453_U275 ( .B1(u4_srl_453_n218), .B2(u4_srl_453_n327), .C1(
        u4_srl_453_n220), .C2(u4_srl_453_n193), .A(u4_srl_453_n328), .ZN(
        u4_srl_453_n326) );
  AOI21_X1 u4_srl_453_U274 ( .B1(u4_srl_453_n325), .B2(u4_srl_453_n326), .A(
        u4_shift_right[8]), .ZN(u4_N5910) );
  AOI22_X1 u4_srl_453_U273 ( .A1(u4_srl_453_n12), .A2(u4_srl_453_n323), .B1(
        u4_srl_453_n14), .B2(u4_srl_453_n324), .ZN(u4_srl_453_n322) );
  OAI221_X1 u4_srl_453_U272 ( .B1(u4_srl_453_n320), .B2(u4_srl_453_n9), .C1(
        u4_srl_453_n321), .C2(u4_srl_453_n8), .A(u4_srl_453_n322), .ZN(
        u4_N5956) );
  AOI22_X1 u4_srl_453_U271 ( .A1(u4_srl_453_n12), .A2(u4_srl_453_n318), .B1(
        u4_srl_453_n14), .B2(u4_srl_453_n319), .ZN(u4_srl_453_n317) );
  OAI221_X1 u4_srl_453_U270 ( .B1(u4_srl_453_n315), .B2(u4_srl_453_n9), .C1(
        u4_srl_453_n316), .C2(u4_srl_453_n8), .A(u4_srl_453_n317), .ZN(
        u4_N5957) );
  AOI22_X1 u4_srl_453_U269 ( .A1(u4_srl_453_n12), .A2(u4_srl_453_n313), .B1(
        u4_srl_453_n14), .B2(u4_srl_453_n314), .ZN(u4_srl_453_n311) );
  OAI221_X1 u4_srl_453_U268 ( .B1(u4_srl_453_n309), .B2(u4_srl_453_n9), .C1(
        u4_srl_453_n310), .C2(u4_srl_453_n8), .A(u4_srl_453_n311), .ZN(
        u4_N5958) );
  INV_X1 u4_srl_453_U267 ( .A(u4_srl_453_n308), .ZN(u4_srl_453_n291) );
  OAI222_X1 u4_srl_453_U266 ( .A1(u4_srl_453_n289), .A2(u4_srl_453_n181), .B1(
        u4_srl_453_n291), .B2(u4_srl_453_n9), .C1(u4_srl_453_n208), .C2(
        u4_srl_453_n299), .ZN(u4_N5959) );
  INV_X1 u4_srl_453_U265 ( .A(u4_srl_453_n307), .ZN(u4_srl_453_n262) );
  INV_X1 u4_srl_453_U264 ( .A(u4_srl_453_n306), .ZN(u4_srl_453_n207) );
  OAI222_X1 u4_srl_453_U263 ( .A1(u4_srl_453_n260), .A2(u4_srl_453_n181), .B1(
        u4_srl_453_n262), .B2(u4_srl_453_n10), .C1(u4_srl_453_n207), .C2(
        u4_srl_453_n299), .ZN(u4_N5960) );
  INV_X1 u4_srl_453_U262 ( .A(u4_srl_453_n305), .ZN(u4_srl_453_n246) );
  INV_X1 u4_srl_453_U261 ( .A(u4_srl_453_n304), .ZN(u4_srl_453_n206) );
  OAI222_X1 u4_srl_453_U260 ( .A1(u4_srl_453_n229), .A2(u4_srl_453_n181), .B1(
        u4_srl_453_n246), .B2(u4_srl_453_n10), .C1(u4_srl_453_n206), .C2(
        u4_srl_453_n299), .ZN(u4_N5961) );
  INV_X1 u4_srl_453_U259 ( .A(u4_srl_453_n303), .ZN(u4_srl_453_n243) );
  INV_X1 u4_srl_453_U258 ( .A(u4_srl_453_n302), .ZN(u4_srl_453_n205) );
  OAI222_X1 u4_srl_453_U257 ( .A1(u4_srl_453_n201), .A2(u4_srl_453_n181), .B1(
        u4_srl_453_n243), .B2(u4_srl_453_n9), .C1(u4_srl_453_n205), .C2(
        u4_srl_453_n299), .ZN(u4_N5962) );
  INV_X1 u4_srl_453_U256 ( .A(u4_srl_453_n301), .ZN(u4_srl_453_n237) );
  INV_X1 u4_srl_453_U255 ( .A(u4_srl_453_n300), .ZN(u4_srl_453_n203) );
  OAI222_X1 u4_srl_453_U254 ( .A1(u4_srl_453_n176), .A2(u4_srl_453_n181), .B1(
        u4_srl_453_n237), .B2(u4_srl_453_n9), .C1(u4_srl_453_n203), .C2(
        u4_srl_453_n299), .ZN(u4_N5963) );
  OAI222_X1 u4_srl_453_U253 ( .A1(u4_srl_453_n297), .A2(u4_srl_453_n10), .B1(
        u4_srl_453_n190), .B2(u4_srl_453_n4), .C1(u4_srl_453_n298), .C2(
        u4_srl_453_n8), .ZN(u4_N5964) );
  OAI222_X1 u4_srl_453_U252 ( .A1(u4_srl_453_n295), .A2(u4_srl_453_n9), .B1(
        u4_srl_453_n189), .B2(u4_srl_453_n4), .C1(u4_srl_453_n296), .C2(
        u4_srl_453_n8), .ZN(u4_N5965) );
  OAI222_X1 u4_srl_453_U251 ( .A1(u4_srl_453_n291), .A2(u4_srl_453_n238), .B1(
        u4_srl_453_n292), .B2(u4_srl_453_n293), .C1(u4_srl_453_n294), .C2(
        u4_srl_453_n242), .ZN(u4_srl_453_n267) );
  OAI22_X1 u4_srl_453_U250 ( .A1(u4_srl_453_n289), .A2(u4_srl_453_n177), .B1(
        u4_srl_453_n290), .B2(u4_srl_453_n179), .ZN(u4_srl_453_n288) );
  AOI221_X1 u4_srl_453_U249 ( .B1(u4_srl_453_n171), .B2(u4_srl_453_n287), .C1(
        u4_srl_453_n267), .C2(u4_srl_453_n174), .A(u4_srl_453_n288), .ZN(
        u4_srl_453_n281) );
  AOI22_X1 u4_srl_453_U248 ( .A1(u4_srl_453_n286), .A2(u4_srl_453_n164), .B1(
        u4_srl_453_n165), .B2(u4_srl_453_n162), .ZN(u4_srl_453_n285) );
  INV_X1 u4_srl_453_U247 ( .A(u4_srl_453_n285), .ZN(u4_srl_453_n284) );
  AOI221_X1 u4_srl_453_U246 ( .B1(u4_srl_453_n218), .B2(u4_srl_453_n283), .C1(
        u4_srl_453_n220), .C2(u4_srl_453_n163), .A(u4_srl_453_n284), .ZN(
        u4_srl_453_n282) );
  AOI21_X1 u4_srl_453_U245 ( .B1(u4_srl_453_n281), .B2(u4_srl_453_n282), .A(
        u4_shift_right[8]), .ZN(u4_N5911) );
  OAI222_X1 u4_srl_453_U244 ( .A1(u4_srl_453_n279), .A2(u4_srl_453_n9), .B1(
        u4_srl_453_n188), .B2(u4_srl_453_n4), .C1(u4_srl_453_n280), .C2(
        u4_srl_453_n8), .ZN(u4_N5966) );
  OAI222_X1 u4_srl_453_U243 ( .A1(u4_srl_453_n277), .A2(u4_srl_453_n9), .B1(
        u4_srl_453_n187), .B2(u4_srl_453_n4), .C1(u4_srl_453_n278), .C2(
        u4_srl_453_n8), .ZN(u4_N5967) );
  OAI222_X1 u4_srl_453_U242 ( .A1(u4_srl_453_n275), .A2(u4_srl_453_n9), .B1(
        u4_srl_453_n186), .B2(u4_srl_453_n4), .C1(u4_srl_453_n276), .C2(
        u4_srl_453_n181), .ZN(u4_N5968) );
  OAI222_X1 u4_srl_453_U241 ( .A1(u4_srl_453_n273), .A2(u4_srl_453_n9), .B1(
        u4_srl_453_n185), .B2(u4_srl_453_n4), .C1(u4_srl_453_n274), .C2(
        u4_srl_453_n181), .ZN(u4_N5969) );
  INV_X1 u4_srl_453_U240 ( .A(u4_srl_453_n210), .ZN(u4_srl_453_n212) );
  NOR2_X1 u4_srl_453_U239 ( .A1(u4_srl_453_n272), .A2(u4_srl_453_n212), .ZN(
        u4_N5970) );
  NOR2_X1 u4_srl_453_U238 ( .A1(u4_srl_453_n271), .A2(u4_srl_453_n212), .ZN(
        u4_N5971) );
  NOR2_X1 u4_srl_453_U237 ( .A1(u4_srl_453_n270), .A2(u4_srl_453_n212), .ZN(
        u4_N5972) );
  NOR2_X1 u4_srl_453_U236 ( .A1(u4_srl_453_n269), .A2(u4_srl_453_n212), .ZN(
        u4_N5973) );
  AND2_X1 u4_srl_453_U235 ( .A1(u4_srl_453_n268), .A2(u4_srl_453_n210), .ZN(
        u4_N5974) );
  AND2_X1 u4_srl_453_U234 ( .A1(u4_srl_453_n267), .A2(u4_srl_453_n210), .ZN(
        u4_N5975) );
  OR2_X1 u4_srl_453_U233 ( .A1(u4_srl_453_n265), .A2(u4_srl_453_n266), .ZN(
        u4_srl_453_n239) );
  OAI222_X1 u4_srl_453_U232 ( .A1(u4_srl_453_n262), .A2(u4_srl_453_n238), .B1(
        u4_srl_453_n263), .B2(u4_srl_453_n239), .C1(u4_srl_453_n264), .C2(
        u4_srl_453_n242), .ZN(u4_srl_453_n249) );
  OAI22_X1 u4_srl_453_U231 ( .A1(u4_srl_453_n260), .A2(u4_srl_453_n177), .B1(
        u4_srl_453_n261), .B2(u4_srl_453_n179), .ZN(u4_srl_453_n259) );
  AOI221_X1 u4_srl_453_U230 ( .B1(u4_srl_453_n171), .B2(u4_srl_453_n258), .C1(
        u4_srl_453_n249), .C2(u4_srl_453_n174), .A(u4_srl_453_n259), .ZN(
        u4_srl_453_n250) );
  AOI22_X1 u4_srl_453_U229 ( .A1(u4_srl_453_n256), .A2(u4_srl_453_n164), .B1(
        u4_srl_453_n257), .B2(u4_srl_453_n162), .ZN(u4_srl_453_n255) );
  INV_X1 u4_srl_453_U228 ( .A(u4_srl_453_n255), .ZN(u4_srl_453_n254) );
  AOI221_X1 u4_srl_453_U227 ( .B1(u4_srl_453_n218), .B2(u4_srl_453_n252), .C1(
        u4_srl_453_n220), .C2(u4_srl_453_n253), .A(u4_srl_453_n254), .ZN(
        u4_srl_453_n251) );
  AOI21_X1 u4_srl_453_U226 ( .B1(u4_srl_453_n250), .B2(u4_srl_453_n251), .A(
        u4_shift_right[8]), .ZN(u4_N5912) );
  AND2_X1 u4_srl_453_U225 ( .A1(u4_srl_453_n249), .A2(u4_srl_453_n210), .ZN(
        u4_N5976) );
  OAI222_X1 u4_srl_453_U224 ( .A1(u4_srl_453_n246), .A2(u4_srl_453_n238), .B1(
        u4_srl_453_n247), .B2(u4_srl_453_n239), .C1(u4_srl_453_n248), .C2(
        u4_srl_453_n242), .ZN(u4_srl_453_n227) );
  AND2_X1 u4_srl_453_U223 ( .A1(u4_srl_453_n227), .A2(u4_srl_453_n210), .ZN(
        u4_N5977) );
  OAI222_X1 u4_srl_453_U222 ( .A1(u4_srl_453_n243), .A2(u4_srl_453_n238), .B1(
        u4_srl_453_n244), .B2(u4_srl_453_n239), .C1(u4_srl_453_n245), .C2(
        u4_srl_453_n242), .ZN(u4_srl_453_n199) );
  AND2_X1 u4_srl_453_U221 ( .A1(u4_srl_453_n199), .A2(u4_srl_453_n210), .ZN(
        u4_N5978) );
  OAI222_X1 u4_srl_453_U220 ( .A1(u4_srl_453_n237), .A2(u4_srl_453_n238), .B1(
        u4_srl_453_n239), .B2(u4_srl_453_n240), .C1(u4_srl_453_n241), .C2(
        u4_srl_453_n242), .ZN(u4_srl_453_n173) );
  AND2_X1 u4_srl_453_U219 ( .A1(u4_srl_453_n173), .A2(u4_srl_453_n210), .ZN(
        u4_N5979) );
  AND2_X1 u4_srl_453_U218 ( .A1(u4_srl_453_n236), .A2(u4_srl_453_n210), .ZN(
        u4_N5980) );
  AND2_X1 u4_srl_453_U217 ( .A1(u4_srl_453_n235), .A2(u4_srl_453_n210), .ZN(
        u4_N5981) );
  AND2_X1 u4_srl_453_U216 ( .A1(u4_srl_453_n234), .A2(u4_srl_453_n210), .ZN(
        u4_N5982) );
  AND2_X1 u4_srl_453_U215 ( .A1(u4_srl_453_n233), .A2(u4_srl_453_n210), .ZN(
        u4_N5983) );
  AND2_X1 u4_srl_453_U214 ( .A1(u4_srl_453_n232), .A2(u4_srl_453_n210), .ZN(
        u4_N5984) );
  AND2_X1 u4_srl_453_U213 ( .A1(u4_srl_453_n231), .A2(u4_srl_453_n210), .ZN(
        u4_N5985) );
  OAI22_X1 u4_srl_453_U212 ( .A1(u4_srl_453_n229), .A2(u4_srl_453_n177), .B1(
        u4_srl_453_n230), .B2(u4_srl_453_n179), .ZN(u4_srl_453_n228) );
  AOI221_X1 u4_srl_453_U211 ( .B1(u4_srl_453_n171), .B2(u4_srl_453_n226), .C1(
        u4_srl_453_n227), .C2(u4_srl_453_n174), .A(u4_srl_453_n228), .ZN(
        u4_srl_453_n216) );
  AOI22_X1 u4_srl_453_U210 ( .A1(u4_srl_453_n224), .A2(u4_srl_453_n164), .B1(
        u4_srl_453_n225), .B2(u4_srl_453_n162), .ZN(u4_srl_453_n223) );
  INV_X1 u4_srl_453_U209 ( .A(u4_srl_453_n223), .ZN(u4_srl_453_n222) );
  AOI221_X1 u4_srl_453_U208 ( .B1(u4_srl_453_n218), .B2(u4_srl_453_n219), .C1(
        u4_srl_453_n220), .C2(u4_srl_453_n221), .A(u4_srl_453_n222), .ZN(
        u4_srl_453_n217) );
  AOI21_X1 u4_srl_453_U207 ( .B1(u4_srl_453_n216), .B2(u4_srl_453_n217), .A(
        u4_shift_right[8]), .ZN(u4_N5913) );
  NOR2_X1 u4_srl_453_U206 ( .A1(u4_srl_453_n215), .A2(u4_srl_453_n212), .ZN(
        u4_N5986) );
  NOR2_X1 u4_srl_453_U205 ( .A1(u4_srl_453_n214), .A2(u4_srl_453_n212), .ZN(
        u4_N5987) );
  NOR2_X1 u4_srl_453_U204 ( .A1(u4_srl_453_n213), .A2(u4_srl_453_n212), .ZN(
        u4_N5988) );
  NOR2_X1 u4_srl_453_U203 ( .A1(u4_srl_453_n211), .A2(u4_srl_453_n212), .ZN(
        u4_N5989) );
  AND2_X1 u4_srl_453_U202 ( .A1(u4_srl_453_n209), .A2(u4_srl_453_n210), .ZN(
        u4_N5990) );
  NOR2_X1 u4_srl_453_U201 ( .A1(u4_srl_453_n208), .A2(u4_srl_453_n204), .ZN(
        u4_N5991) );
  NOR2_X1 u4_srl_453_U200 ( .A1(u4_srl_453_n207), .A2(u4_srl_453_n204), .ZN(
        u4_N5992) );
  NOR2_X1 u4_srl_453_U199 ( .A1(u4_srl_453_n206), .A2(u4_srl_453_n204), .ZN(
        u4_N5993) );
  NOR2_X1 u4_srl_453_U198 ( .A1(u4_srl_453_n205), .A2(u4_srl_453_n204), .ZN(
        u4_N5994) );
  NOR2_X1 u4_srl_453_U197 ( .A1(u4_srl_453_n203), .A2(u4_srl_453_n204), .ZN(
        u4_N5995) );
  OAI22_X1 u4_srl_453_U196 ( .A1(u4_srl_453_n201), .A2(u4_srl_453_n177), .B1(
        u4_srl_453_n202), .B2(u4_srl_453_n179), .ZN(u4_srl_453_n200) );
  AOI221_X1 u4_srl_453_U195 ( .B1(u4_srl_453_n171), .B2(u4_srl_453_n198), .C1(
        u4_srl_453_n199), .C2(u4_srl_453_n174), .A(u4_srl_453_n200), .ZN(
        u4_srl_453_n191) );
  OAI22_X1 u4_srl_453_U194 ( .A1(u4_srl_453_n196), .A2(u4_srl_453_n168), .B1(
        u4_srl_453_n197), .B2(u4_srl_453_n170), .ZN(u4_srl_453_n195) );
  AOI221_X1 u4_srl_453_U193 ( .B1(u4_srl_453_n162), .B2(u4_srl_453_n193), .C1(
        u4_srl_453_n164), .C2(u4_srl_453_n194), .A(u4_srl_453_n195), .ZN(
        u4_srl_453_n192) );
  AOI21_X1 u4_srl_453_U192 ( .B1(u4_srl_453_n191), .B2(u4_srl_453_n192), .A(
        u4_shift_right[8]), .ZN(u4_N5914) );
  NOR2_X1 u4_srl_453_U191 ( .A1(u4_srl_453_n190), .A2(u4_srl_453_n8), .ZN(
        u4_N5996) );
  NOR2_X1 u4_srl_453_U190 ( .A1(u4_srl_453_n189), .A2(u4_srl_453_n8), .ZN(
        u4_N5997) );
  NOR2_X1 u4_srl_453_U189 ( .A1(u4_srl_453_n188), .A2(u4_srl_453_n8), .ZN(
        u4_N5998) );
  NOR2_X1 u4_srl_453_U188 ( .A1(u4_srl_453_n187), .A2(u4_srl_453_n8), .ZN(
        u4_N5999) );
  NOR2_X1 u4_srl_453_U187 ( .A1(u4_srl_453_n186), .A2(u4_srl_453_n8), .ZN(
        u4_N6000) );
  NOR2_X1 u4_srl_453_U186 ( .A1(u4_srl_453_n185), .A2(u4_srl_453_n8), .ZN(
        u4_N6001) );
  NOR2_X1 u4_srl_453_U185 ( .A1(u4_srl_453_n184), .A2(u4_srl_453_n8), .ZN(
        u4_N6002) );
  NOR2_X1 u4_srl_453_U184 ( .A1(u4_srl_453_n183), .A2(u4_srl_453_n8), .ZN(
        u4_N6003) );
  NOR2_X1 u4_srl_453_U183 ( .A1(u4_srl_453_n182), .A2(u4_srl_453_n8), .ZN(
        u4_N6004) );
  NOR2_X1 u4_srl_453_U182 ( .A1(u4_srl_453_n180), .A2(u4_srl_453_n8), .ZN(
        u4_N6005) );
  OAI22_X1 u4_srl_453_U181 ( .A1(u4_srl_453_n176), .A2(u4_srl_453_n177), .B1(
        u4_srl_453_n178), .B2(u4_srl_453_n179), .ZN(u4_srl_453_n175) );
  AOI221_X1 u4_srl_453_U180 ( .B1(u4_srl_453_n171), .B2(u4_srl_453_n172), .C1(
        u4_srl_453_n173), .C2(u4_srl_453_n174), .A(u4_srl_453_n175), .ZN(
        u4_srl_453_n160) );
  OAI22_X1 u4_srl_453_U179 ( .A1(u4_srl_453_n167), .A2(u4_srl_453_n168), .B1(
        u4_srl_453_n169), .B2(u4_srl_453_n170), .ZN(u4_srl_453_n166) );
  AOI221_X1 u4_srl_453_U178 ( .B1(u4_srl_453_n162), .B2(u4_srl_453_n163), .C1(
        u4_srl_453_n164), .C2(u4_srl_453_n165), .A(u4_srl_453_n166), .ZN(
        u4_srl_453_n161) );
  AOI21_X1 u4_srl_453_U177 ( .B1(u4_srl_453_n160), .B2(u4_srl_453_n161), .A(
        u4_shift_right[8]), .ZN(u4_N5915) );
  INV_X4 u4_srl_453_U176 ( .A(n6445), .ZN(u4_srl_453_n159) );
  INV_X4 u4_srl_453_U175 ( .A(n6444), .ZN(u4_srl_453_n158) );
  INV_X4 u4_srl_453_U174 ( .A(n6443), .ZN(u4_srl_453_n157) );
  INV_X4 u4_srl_453_U173 ( .A(n6442), .ZN(u4_srl_453_n156) );
  INV_X4 u4_srl_453_U172 ( .A(n6441), .ZN(u4_srl_453_n155) );
  INV_X4 u4_srl_453_U171 ( .A(n6440), .ZN(u4_srl_453_n154) );
  INV_X4 u4_srl_453_U170 ( .A(n6439), .ZN(u4_srl_453_n153) );
  INV_X4 u4_srl_453_U169 ( .A(n6438), .ZN(u4_srl_453_n152) );
  INV_X4 u4_srl_453_U168 ( .A(n6437), .ZN(u4_srl_453_n151) );
  INV_X4 u4_srl_453_U167 ( .A(n6436), .ZN(u4_srl_453_n150) );
  INV_X4 u4_srl_453_U166 ( .A(n6435), .ZN(u4_srl_453_n149) );
  INV_X4 u4_srl_453_U165 ( .A(n6434), .ZN(u4_srl_453_n148) );
  INV_X4 u4_srl_453_U164 ( .A(n6433), .ZN(u4_srl_453_n147) );
  INV_X4 u4_srl_453_U163 ( .A(n6432), .ZN(u4_srl_453_n146) );
  INV_X4 u4_srl_453_U162 ( .A(n6431), .ZN(u4_srl_453_n145) );
  INV_X4 u4_srl_453_U161 ( .A(n6430), .ZN(u4_srl_453_n144) );
  INV_X4 u4_srl_453_U160 ( .A(n6429), .ZN(u4_srl_453_n143) );
  INV_X4 u4_srl_453_U159 ( .A(n6428), .ZN(u4_srl_453_n142) );
  INV_X4 u4_srl_453_U158 ( .A(n6427), .ZN(u4_srl_453_n141) );
  INV_X4 u4_srl_453_U157 ( .A(n6426), .ZN(u4_srl_453_n140) );
  INV_X4 u4_srl_453_U156 ( .A(n6425), .ZN(u4_srl_453_n139) );
  INV_X4 u4_srl_453_U155 ( .A(n6424), .ZN(u4_srl_453_n138) );
  INV_X4 u4_srl_453_U154 ( .A(n6423), .ZN(u4_srl_453_n137) );
  INV_X4 u4_srl_453_U153 ( .A(n6422), .ZN(u4_srl_453_n136) );
  INV_X4 u4_srl_453_U152 ( .A(n6421), .ZN(u4_srl_453_n135) );
  INV_X4 u4_srl_453_U151 ( .A(n6419), .ZN(u4_srl_453_n134) );
  INV_X4 u4_srl_453_U150 ( .A(n6418), .ZN(u4_srl_453_n133) );
  INV_X4 u4_srl_453_U149 ( .A(n6417), .ZN(u4_srl_453_n132) );
  INV_X4 u4_srl_453_U148 ( .A(n6416), .ZN(u4_srl_453_n131) );
  INV_X4 u4_srl_453_U147 ( .A(n6415), .ZN(u4_srl_453_n130) );
  INV_X4 u4_srl_453_U146 ( .A(n6414), .ZN(u4_srl_453_n129) );
  INV_X4 u4_srl_453_U145 ( .A(n6413), .ZN(u4_srl_453_n128) );
  INV_X4 u4_srl_453_U144 ( .A(n6411), .ZN(u4_srl_453_n127) );
  INV_X4 u4_srl_453_U143 ( .A(n6410), .ZN(u4_srl_453_n126) );
  INV_X4 u4_srl_453_U142 ( .A(n6409), .ZN(u4_srl_453_n125) );
  INV_X4 u4_srl_453_U141 ( .A(n6408), .ZN(u4_srl_453_n124) );
  INV_X4 u4_srl_453_U140 ( .A(n6407), .ZN(u4_srl_453_n123) );
  INV_X4 u4_srl_453_U139 ( .A(n6406), .ZN(u4_srl_453_n122) );
  INV_X4 u4_srl_453_U138 ( .A(n6405), .ZN(u4_srl_453_n121) );
  INV_X4 u4_srl_453_U137 ( .A(fract_denorm[50]), .ZN(u4_srl_453_n120) );
  INV_X4 u4_srl_453_U136 ( .A(fract_denorm[51]), .ZN(u4_srl_453_n119) );
  INV_X4 u4_srl_453_U135 ( .A(fract_denorm[74]), .ZN(u4_srl_453_n118) );
  INV_X4 u4_srl_453_U134 ( .A(fract_denorm[82]), .ZN(u4_srl_453_n117) );
  INV_X4 u4_srl_453_U133 ( .A(fract_denorm[66]), .ZN(u4_srl_453_n116) );
  INV_X4 u4_srl_453_U132 ( .A(fract_denorm[58]), .ZN(u4_srl_453_n115) );
  INV_X4 u4_srl_453_U131 ( .A(fract_denorm[52]), .ZN(u4_srl_453_n114) );
  INV_X4 u4_srl_453_U130 ( .A(fract_denorm[71]), .ZN(u4_srl_453_n113) );
  INV_X4 u4_srl_453_U129 ( .A(fract_denorm[73]), .ZN(u4_srl_453_n112) );
  INV_X4 u4_srl_453_U128 ( .A(fract_denorm[72]), .ZN(u4_srl_453_n111) );
  INV_X4 u4_srl_453_U127 ( .A(fract_denorm[70]), .ZN(u4_srl_453_n110) );
  INV_X4 u4_srl_453_U126 ( .A(fract_denorm[69]), .ZN(u4_srl_453_n109) );
  INV_X4 u4_srl_453_U125 ( .A(fract_denorm[68]), .ZN(u4_srl_453_n108) );
  INV_X4 u4_srl_453_U124 ( .A(fract_denorm[67]), .ZN(u4_srl_453_n107) );
  INV_X4 u4_srl_453_U123 ( .A(fract_denorm[63]), .ZN(u4_srl_453_n106) );
  INV_X4 u4_srl_453_U122 ( .A(fract_denorm[65]), .ZN(u4_srl_453_n105) );
  INV_X4 u4_srl_453_U121 ( .A(fract_denorm[64]), .ZN(u4_srl_453_n104) );
  INV_X4 u4_srl_453_U120 ( .A(fract_denorm[62]), .ZN(u4_srl_453_n103) );
  INV_X4 u4_srl_453_U119 ( .A(fract_denorm[61]), .ZN(u4_srl_453_n102) );
  INV_X4 u4_srl_453_U118 ( .A(fract_denorm[60]), .ZN(u4_srl_453_n101) );
  INV_X4 u4_srl_453_U117 ( .A(fract_denorm[59]), .ZN(u4_srl_453_n100) );
  INV_X4 u4_srl_453_U116 ( .A(fract_denorm[79]), .ZN(u4_srl_453_n99) );
  INV_X4 u4_srl_453_U115 ( .A(fract_denorm[81]), .ZN(u4_srl_453_n98) );
  INV_X4 u4_srl_453_U114 ( .A(fract_denorm[80]), .ZN(u4_srl_453_n97) );
  INV_X4 u4_srl_453_U113 ( .A(fract_denorm[78]), .ZN(u4_srl_453_n96) );
  INV_X4 u4_srl_453_U112 ( .A(fract_denorm[77]), .ZN(u4_srl_453_n95) );
  INV_X4 u4_srl_453_U111 ( .A(fract_denorm[76]), .ZN(u4_srl_453_n94) );
  INV_X4 u4_srl_453_U110 ( .A(fract_denorm[75]), .ZN(u4_srl_453_n93) );
  INV_X4 u4_srl_453_U109 ( .A(fract_denorm[87]), .ZN(u4_srl_453_n92) );
  INV_X4 u4_srl_453_U108 ( .A(fract_denorm[89]), .ZN(u4_srl_453_n91) );
  INV_X4 u4_srl_453_U107 ( .A(fract_denorm[88]), .ZN(u4_srl_453_n90) );
  INV_X4 u4_srl_453_U106 ( .A(fract_denorm[86]), .ZN(u4_srl_453_n89) );
  INV_X4 u4_srl_453_U105 ( .A(fract_denorm[85]), .ZN(u4_srl_453_n88) );
  INV_X4 u4_srl_453_U104 ( .A(fract_denorm[84]), .ZN(u4_srl_453_n87) );
  INV_X4 u4_srl_453_U103 ( .A(fract_denorm[83]), .ZN(u4_srl_453_n86) );
  INV_X4 u4_srl_453_U102 ( .A(fract_denorm[55]), .ZN(u4_srl_453_n85) );
  INV_X4 u4_srl_453_U101 ( .A(fract_denorm[57]), .ZN(u4_srl_453_n84) );
  INV_X4 u4_srl_453_U100 ( .A(fract_denorm[56]), .ZN(u4_srl_453_n83) );
  INV_X4 u4_srl_453_U99 ( .A(fract_denorm[54]), .ZN(u4_srl_453_n82) );
  INV_X4 u4_srl_453_U98 ( .A(fract_denorm[53]), .ZN(u4_srl_453_n81) );
  INV_X4 u4_srl_453_U97 ( .A(n6367), .ZN(u4_srl_453_n80) );
  INV_X4 u4_srl_453_U96 ( .A(fract_denorm[98]), .ZN(u4_srl_453_n79) );
  INV_X4 u4_srl_453_U95 ( .A(fract_denorm[100]), .ZN(u4_srl_453_n78) );
  INV_X4 u4_srl_453_U94 ( .A(fract_denorm[102]), .ZN(u4_srl_453_n77) );
  INV_X4 u4_srl_453_U93 ( .A(fract_denorm[101]), .ZN(u4_srl_453_n76) );
  INV_X4 u4_srl_453_U92 ( .A(fract_denorm[99]), .ZN(u4_srl_453_n75) );
  INV_X4 u4_srl_453_U91 ( .A(fract_denorm[90]), .ZN(u4_srl_453_n74) );
  INV_X4 u4_srl_453_U90 ( .A(fract_denorm[95]), .ZN(u4_srl_453_n73) );
  INV_X4 u4_srl_453_U89 ( .A(fract_denorm[97]), .ZN(u4_srl_453_n72) );
  INV_X4 u4_srl_453_U88 ( .A(fract_denorm[96]), .ZN(u4_srl_453_n71) );
  INV_X4 u4_srl_453_U87 ( .A(fract_denorm[94]), .ZN(u4_srl_453_n70) );
  INV_X4 u4_srl_453_U86 ( .A(fract_denorm[93]), .ZN(u4_srl_453_n69) );
  INV_X4 u4_srl_453_U85 ( .A(fract_denorm[92]), .ZN(u4_srl_453_n68) );
  INV_X4 u4_srl_453_U84 ( .A(fract_denorm[91]), .ZN(u4_srl_453_n67) );
  INV_X4 u4_srl_453_U83 ( .A(n6351), .ZN(u4_srl_453_n66) );
  INV_X4 u4_srl_453_U82 ( .A(n6350), .ZN(u4_srl_453_n65) );
  INV_X4 u4_srl_453_U81 ( .A(n6349), .ZN(u4_srl_453_n64) );
  INV_X4 u4_srl_453_U80 ( .A(n6348), .ZN(u4_srl_453_n63) );
  INV_X4 u4_srl_453_U79 ( .A(n6347), .ZN(u4_srl_453_n62) );
  INV_X4 u4_srl_453_U78 ( .A(n6346), .ZN(u4_srl_453_n61) );
  INV_X4 u4_srl_453_U77 ( .A(n6345), .ZN(u4_srl_453_n60) );
  INV_X4 u4_srl_453_U76 ( .A(u4_srl_453_n376), .ZN(u4_srl_453_n383) );
  INV_X4 u4_srl_453_U75 ( .A(u4_srl_453_n859), .ZN(u4_srl_453_n174) );
  AND2_X4 u4_srl_453_U74 ( .A1(u4_srl_453_n16), .A2(u4_srl_453_n794), .ZN(
        u4_srl_453_n162) );
  AND2_X4 u4_srl_453_U73 ( .A1(u4_srl_453_n409), .A2(u4_srl_453_n794), .ZN(
        u4_srl_453_n164) );
  INV_X4 u4_srl_453_U72 ( .A(u4_srl_453_n4), .ZN(u4_srl_453_n14) );
  INV_X4 u4_srl_453_U71 ( .A(u4_srl_453_n409), .ZN(u4_srl_453_n59) );
  INV_X4 u4_srl_453_U70 ( .A(u4_srl_453_n5), .ZN(u4_srl_453_n9) );
  INV_X4 u4_srl_453_U69 ( .A(u4_srl_453_n5), .ZN(u4_srl_453_n10) );
  INV_X4 u4_srl_453_U68 ( .A(u4_srl_453_n11), .ZN(u4_srl_453_n12) );
  INV_X4 u4_srl_453_U67 ( .A(u4_srl_453_n41), .ZN(u4_srl_453_n39) );
  INV_X4 u4_srl_453_U66 ( .A(u4_srl_453_n41), .ZN(u4_srl_453_n37) );
  INV_X4 u4_srl_453_U65 ( .A(u4_srl_453_n41), .ZN(u4_srl_453_n40) );
  INV_X4 u4_srl_453_U64 ( .A(u4_srl_453_n3), .ZN(u4_srl_453_n26) );
  INV_X4 u4_srl_453_U63 ( .A(u4_srl_453_n3), .ZN(u4_srl_453_n27) );
  INV_X4 u4_srl_453_U62 ( .A(u4_srl_453_n3), .ZN(u4_srl_453_n28) );
  INV_X4 u4_srl_453_U61 ( .A(u4_srl_453_n24), .ZN(u4_srl_453_n20) );
  INV_X4 u4_srl_453_U60 ( .A(u4_srl_453_n24), .ZN(u4_srl_453_n22) );
  INV_X4 u4_srl_453_U59 ( .A(u4_srl_453_n24), .ZN(u4_srl_453_n23) );
  INV_X4 u4_srl_453_U58 ( .A(u4_srl_453_n18), .ZN(u4_srl_453_n16) );
  INV_X4 u4_srl_453_U57 ( .A(u4_srl_453_n312), .ZN(u4_srl_453_n11) );
  INV_X4 u4_srl_453_U56 ( .A(u4_srl_453_n4), .ZN(u4_srl_453_n13) );
  INV_X4 u4_srl_453_U55 ( .A(u4_srl_453_n3), .ZN(u4_srl_453_n25) );
  INV_X4 u4_srl_453_U54 ( .A(u4_srl_453_n58), .ZN(u4_srl_453_n57) );
  INV_X4 u4_srl_453_U53 ( .A(u4_srl_453_n6), .ZN(u4_srl_453_n41) );
  INV_X4 u4_srl_453_U52 ( .A(u4_srl_453_n393), .ZN(u4_srl_453_n18) );
  INV_X4 u4_srl_453_U51 ( .A(u4_srl_453_n24), .ZN(u4_srl_453_n21) );
  INV_X4 u4_srl_453_U50 ( .A(u4_srl_453_n1), .ZN(u4_srl_453_n42) );
  INV_X4 u4_srl_453_U49 ( .A(u4_srl_453_n41), .ZN(u4_srl_453_n38) );
  INV_X4 u4_srl_453_U48 ( .A(u4_srl_453_n394), .ZN(u4_srl_453_n24) );
  INV_X4 u4_srl_453_U47 ( .A(u4_srl_453_n1), .ZN(u4_srl_453_n43) );
  INV_X4 u4_srl_453_U46 ( .A(u4_srl_453_n1), .ZN(u4_srl_453_n46) );
  INV_X4 u4_srl_453_U45 ( .A(u4_srl_453_n58), .ZN(u4_srl_453_n56) );
  INV_X4 u4_srl_453_U44 ( .A(u4_srl_453_n409), .ZN(u4_srl_453_n58) );
  INV_X4 u4_srl_453_U43 ( .A(u4_srl_453_n393), .ZN(u4_srl_453_n19) );
  INV_X4 u4_srl_453_U42 ( .A(u4_srl_453_n7), .ZN(u4_srl_453_n8) );
  INV_X4 u4_srl_453_U41 ( .A(u4_srl_453_n55), .ZN(u4_srl_453_n51) );
  INV_X4 u4_srl_453_U40 ( .A(u4_srl_453_n55), .ZN(u4_srl_453_n52) );
  INV_X4 u4_srl_453_U39 ( .A(u4_srl_453_n1), .ZN(u4_srl_453_n45) );
  INV_X4 u4_srl_453_U38 ( .A(u4_srl_453_n18), .ZN(u4_srl_453_n17) );
  INV_X4 u4_srl_453_U37 ( .A(u4_srl_453_n19), .ZN(u4_srl_453_n15) );
  INV_X4 u4_srl_453_U36 ( .A(u4_srl_453_n181), .ZN(u4_srl_453_n7) );
  INV_X4 u4_srl_453_U35 ( .A(u4_srl_453_n396), .ZN(u4_srl_453_n54) );
  INV_X4 u4_srl_453_U34 ( .A(u4_srl_453_n1), .ZN(u4_srl_453_n44) );
  NAND2_X2 u4_srl_453_U33 ( .A1(u4_srl_453_n878), .A2(u4_srl_453_n879), .ZN(
        u4_srl_453_n6) );
  NOR2_X2 u4_srl_453_U32 ( .A1(u4_shift_right[0]), .A2(u4_srl_453_n878), .ZN(
        u4_srl_453_n396) );
  INV_X4 u4_srl_453_U31 ( .A(u4_srl_453_n396), .ZN(u4_srl_453_n55) );
  INV_X4 u4_srl_453_U30 ( .A(u4_srl_453_n35), .ZN(u4_srl_453_n29) );
  INV_X4 u4_srl_453_U29 ( .A(u4_srl_453_n34), .ZN(u4_srl_453_n31) );
  INV_X4 u4_srl_453_U28 ( .A(u4_srl_453_n41), .ZN(u4_srl_453_n36) );
  AND2_X4 u4_srl_453_U27 ( .A1(u4_srl_453_n386), .A2(u4_shift_right[4]), .ZN(
        u4_srl_453_n5) );
  INV_X4 u4_srl_453_U26 ( .A(u4_srl_453_n31), .ZN(u4_srl_453_n33) );
  OR2_X4 u4_srl_453_U25 ( .A1(u4_srl_453_n299), .A2(u4_shift_right[4]), .ZN(
        u4_srl_453_n4) );
  OR2_X4 u4_srl_453_U24 ( .A1(u4_shift_right[2]), .A2(u4_srl_453_n833), .ZN(
        u4_srl_453_n3) );
  NAND2_X4 u4_srl_453_U23 ( .A1(u4_srl_453_n878), .A2(u4_shift_right[0]), .ZN(
        u4_srl_453_n2) );
  OR2_X4 u4_srl_453_U22 ( .A1(u4_srl_453_n879), .A2(u4_srl_453_n878), .ZN(
        u4_srl_453_n1) );
  NOR2_X2 u4_srl_453_U21 ( .A1(u4_srl_453_n174), .A2(u4_shift_right[8]), .ZN(
        u4_srl_453_n210) );
  NOR2_X2 u4_srl_453_U20 ( .A1(u4_srl_453_n242), .A2(u4_srl_453_n174), .ZN(
        u4_srl_453_n171) );
  NAND2_X2 u4_srl_453_U19 ( .A1(u4_srl_453_n794), .A2(u4_srl_453_n23), .ZN(
        u4_srl_453_n170) );
  NAND2_X2 u4_srl_453_U18 ( .A1(u4_srl_453_n26), .A2(u4_srl_453_n794), .ZN(
        u4_srl_453_n168) );
  NOR2_X2 u4_srl_453_U17 ( .A1(u4_srl_453_n383), .A2(u4_srl_453_n238), .ZN(
        u4_srl_453_n408) );
  INV_X4 u4_srl_453_U16 ( .A(u4_shift_right[4]), .ZN(u4_srl_453_n392) );
  INV_X4 u4_srl_453_U15 ( .A(u4_srl_453_n53), .ZN(u4_srl_453_n47) );
  INV_X4 u4_srl_453_U14 ( .A(u4_srl_453_n2), .ZN(u4_srl_453_n35) );
  NAND2_X2 u4_srl_453_U13 ( .A1(u4_srl_453_n266), .A2(u4_srl_453_n392), .ZN(
        u4_srl_453_n238) );
  NAND2_X2 u4_srl_453_U12 ( .A1(u4_srl_453_n266), .A2(u4_shift_right[4]), .ZN(
        u4_srl_453_n242) );
  INV_X4 u4_srl_453_U11 ( .A(u4_srl_453_n33), .ZN(u4_srl_453_n32) );
  NAND2_X2 u4_srl_453_U10 ( .A1(u4_srl_453_n801), .A2(u4_shift_right[4]), .ZN(
        u4_srl_453_n177) );
  NAND2_X2 u4_srl_453_U9 ( .A1(u4_srl_453_n801), .A2(u4_srl_453_n392), .ZN(
        u4_srl_453_n179) );
  INV_X4 u4_srl_453_U8 ( .A(u4_srl_453_n34), .ZN(u4_srl_453_n30) );
  INV_X4 u4_srl_453_U7 ( .A(u4_srl_453_n53), .ZN(u4_srl_453_n49) );
  INV_X4 u4_srl_453_U6 ( .A(u4_srl_453_n53), .ZN(u4_srl_453_n48) );
  INV_X4 u4_srl_453_U5 ( .A(u4_srl_453_n54), .ZN(u4_srl_453_n50) );
  INV_X4 u4_srl_453_U4 ( .A(u4_srl_453_n51), .ZN(u4_srl_453_n53) );
  INV_X4 u4_srl_453_U3 ( .A(u4_srl_453_n2), .ZN(u4_srl_453_n34) );
  OR3_X1 u4_sll_482_U88 ( .A1(u4_f2i_shft_8_), .A2(u4_f2i_shft_9_), .A3(
        u4_f2i_shft_7_), .ZN(u4_sll_482_n57) );
  NAND2_X1 u4_sll_482_U87 ( .A1(u4_sll_482_n57), .A2(u4_sll_482_n44), .ZN(
        u4_sll_482_n46) );
  NAND3_X1 u4_sll_482_U86 ( .A1(u4_f2i_shft_8_), .A2(u4_f2i_shft_7_), .A3(
        u4_f2i_shft_9_), .ZN(u4_sll_482_n56) );
  NAND2_X1 u4_sll_482_U85 ( .A1(u4_f2i_shft_10_), .A2(u4_sll_482_n56), .ZN(
        u4_sll_482_n45) );
  NAND2_X1 u4_sll_482_U84 ( .A1(n4349), .A2(u4_sll_482_n45), .ZN(
        u4_sll_482_n55) );
  NAND2_X1 u4_sll_482_U83 ( .A1(u4_sll_482_n46), .A2(u4_sll_482_n55), .ZN(
        u4_sll_482_temp_int_SH_0_) );
  AND2_X1 u4_sll_482_U82 ( .A1(n6446), .A2(u4_sll_482_n11), .ZN(
        u4_sll_482_ML_int_1__0_) );
  AND2_X1 u4_sll_482_U81 ( .A1(fract_denorm[105]), .A2(u4_sll_482_n6), .ZN(
        u4_sll_482_MR_int_1__113_) );
  NAND2_X1 u4_sll_482_U80 ( .A1(u4_f2i_shft_1_), .A2(u4_sll_482_n45), .ZN(
        u4_sll_482_n54) );
  NAND2_X1 u4_sll_482_U79 ( .A1(u4_sll_482_ML_int_1__0_), .A2(u4_sll_482_n1), 
        .ZN(u4_sll_482_n51) );
  NAND2_X1 u4_sll_482_U78 ( .A1(u4_sll_482_ML_int_1__1_), .A2(u4_sll_482_n1), 
        .ZN(u4_sll_482_n50) );
  NAND2_X1 u4_sll_482_U77 ( .A1(u4_f2i_shft_2_), .A2(u4_sll_482_n45), .ZN(
        u4_sll_482_n53) );
  NAND2_X1 u4_sll_482_U76 ( .A1(u4_sll_482_ML_int_2__3_), .A2(u4_sll_482_n2), 
        .ZN(u4_sll_482_n48) );
  NAND2_X1 u4_sll_482_U75 ( .A1(u4_f2i_shft_3_), .A2(u4_sll_482_n45), .ZN(
        u4_sll_482_n52) );
  NAND2_X1 u4_sll_482_U74 ( .A1(u4_sll_482_n46), .A2(u4_sll_482_n52), .ZN(
        u4_sll_482_temp_int_SH_3_) );
  NAND2_X1 u4_sll_482_U73 ( .A1(u4_sll_482_n2), .A2(u4_sll_482_n33), .ZN(
        u4_sll_482_n49) );
  NOR2_X1 u4_sll_482_U72 ( .A1(u4_sll_482_n49), .A2(u4_sll_482_n51), .ZN(
        u4_sll_482_ML_int_4__0_) );
  NOR2_X1 u4_sll_482_U71 ( .A1(u4_sll_482_n49), .A2(u4_sll_482_n50), .ZN(
        u4_sll_482_ML_int_4__1_) );
  NOR2_X1 u4_sll_482_U70 ( .A1(u4_sll_482_n38), .A2(u4_sll_482_n49), .ZN(
        u4_sll_482_ML_int_4__2_) );
  NOR2_X1 u4_sll_482_U69 ( .A1(u4_sll_482_n30), .A2(u4_sll_482_n48), .ZN(
        u4_sll_482_ML_int_4__3_) );
  AND2_X1 u4_sll_482_U68 ( .A1(u4_sll_482_ML_int_3__4_), .A2(u4_sll_482_n33), 
        .ZN(u4_sll_482_ML_int_4__4_) );
  AND2_X1 u4_sll_482_U67 ( .A1(u4_sll_482_ML_int_3__5_), .A2(u4_sll_482_n33), 
        .ZN(u4_sll_482_ML_int_4__5_) );
  NAND2_X1 u4_sll_482_U66 ( .A1(u4_f2i_shft_4_), .A2(u4_sll_482_n45), .ZN(
        u4_sll_482_n47) );
  NAND2_X1 u4_sll_482_U65 ( .A1(u4_sll_482_n46), .A2(u4_sll_482_n47), .ZN(
        u4_sll_482_temp_int_SH_4_) );
  AND2_X1 u4_sll_482_U64 ( .A1(u4_sll_482_ML_int_4__11_), .A2(u4_sll_482_n34), 
        .ZN(u4_sll_482_ML_int_5__11_) );
  AND2_X1 u4_sll_482_U63 ( .A1(u4_sll_482_ML_int_4__12_), .A2(u4_sll_482_n34), 
        .ZN(u4_sll_482_ML_int_5__12_) );
  AND2_X1 u4_sll_482_U62 ( .A1(u4_sll_482_ML_int_4__13_), .A2(u4_sll_482_n34), 
        .ZN(u4_sll_482_ML_int_5__13_) );
  AND2_X1 u4_sll_482_U61 ( .A1(u4_sll_482_ML_int_4__14_), .A2(u4_sll_482_n34), 
        .ZN(u4_sll_482_ML_int_5__14_) );
  AND2_X1 u4_sll_482_U60 ( .A1(u4_sll_482_ML_int_4__15_), .A2(u4_sll_482_n34), 
        .ZN(u4_sll_482_ML_int_5__15_) );
  AND2_X1 u4_sll_482_U59 ( .A1(u4_sll_482_ML_int_7__107_), .A2(u4_sll_482_n44), 
        .ZN(u4_exp_f2i_1[107]) );
  AND2_X1 u4_sll_482_U58 ( .A1(u4_sll_482_ML_int_7__108_), .A2(u4_sll_482_n44), 
        .ZN(u4_exp_f2i_1[108]) );
  AND2_X1 u4_sll_482_U57 ( .A1(u4_sll_482_ML_int_7__109_), .A2(u4_sll_482_n44), 
        .ZN(u4_exp_f2i_1[109]) );
  AND2_X1 u4_sll_482_U56 ( .A1(u4_sll_482_ML_int_7__110_), .A2(u4_sll_482_n44), 
        .ZN(u4_exp_f2i_1[110]) );
  AND2_X1 u4_sll_482_U55 ( .A1(u4_sll_482_ML_int_7__111_), .A2(u4_sll_482_n44), 
        .ZN(u4_exp_f2i_1[111]) );
  AND2_X1 u4_sll_482_U54 ( .A1(u4_sll_482_ML_int_7__112_), .A2(u4_sll_482_n44), 
        .ZN(u4_exp_f2i_1[112]) );
  AND2_X1 u4_sll_482_U53 ( .A1(u4_sll_482_ML_int_7__113_), .A2(u4_sll_482_n44), 
        .ZN(u4_exp_f2i_1[113]) );
  AND2_X1 u4_sll_482_U52 ( .A1(u4_sll_482_ML_int_7__114_), .A2(u4_sll_482_n44), 
        .ZN(u4_exp_f2i_1[114]) );
  AND2_X1 u4_sll_482_U51 ( .A1(u4_sll_482_ML_int_7__115_), .A2(u4_sll_482_n44), 
        .ZN(u4_exp_f2i_1[115]) );
  AND2_X1 u4_sll_482_U50 ( .A1(u4_sll_482_ML_int_7__116_), .A2(u4_sll_482_n44), 
        .ZN(u4_exp_f2i_1[116]) );
  AND2_X1 u4_sll_482_U49 ( .A1(u4_sll_482_ML_int_7__117_), .A2(u4_sll_482_n44), 
        .ZN(u4_exp_f2i_1[117]) );
  OAI21_X1 u4_sll_482_U48 ( .B1(u4_f2i_shft_5_), .B2(u4_sll_482_n43), .A(
        u4_sll_482_n45), .ZN(u4_sll_482_SHMAG[5]) );
  OAI21_X1 u4_sll_482_U47 ( .B1(u4_f2i_shft_6_), .B2(u4_sll_482_n43), .A(
        u4_sll_482_n45), .ZN(u4_sll_482_SHMAG[6]) );
  INV_X4 u4_sll_482_U46 ( .A(u4_f2i_shft_10_), .ZN(u4_sll_482_n44) );
  INV_X4 u4_sll_482_U45 ( .A(u4_sll_482_n46), .ZN(u4_sll_482_n43) );
  INV_X4 u4_sll_482_U44 ( .A(u4_sll_482_SHMAG[6]), .ZN(u4_sll_482_n42) );
  INV_X4 u4_sll_482_U43 ( .A(u4_sll_482_SHMAG[5]), .ZN(u4_sll_482_n41) );
  INV_X4 u4_sll_482_U42 ( .A(u4_sll_482_n48), .ZN(u4_sll_482_n40) );
  INV_X4 u4_sll_482_U41 ( .A(u4_sll_482_n50), .ZN(u4_sll_482_n39) );
  INV_X4 u4_sll_482_U40 ( .A(u4_sll_482_ML_int_2__2_), .ZN(u4_sll_482_n38) );
  INV_X4 u4_sll_482_U39 ( .A(u4_sll_482_n51), .ZN(u4_sll_482_n37) );
  AND2_X4 u4_sll_482_U38 ( .A1(u4_sll_482_n29), .A2(u4_sll_482_ML_int_2__113_), 
        .ZN(u4_sll_482_n5) );
  AND2_X4 u4_sll_482_U37 ( .A1(u4_sll_482_n15), .A2(u4_sll_482_MR_int_1__113_), 
        .ZN(u4_sll_482_n4) );
  INV_X4 u4_sll_482_U36 ( .A(u4_sll_482_n14), .ZN(u4_sll_482_n13) );
  INV_X4 u4_sll_482_U35 ( .A(u4_sll_482_n1), .ZN(u4_sll_482_n21) );
  INV_X4 u4_sll_482_U34 ( .A(u4_sll_482_n1), .ZN(u4_sll_482_n22) );
  INV_X4 u4_sll_482_U33 ( .A(u4_sll_482_n34), .ZN(u4_sll_482_n36) );
  INV_X4 u4_sll_482_U32 ( .A(u4_sll_482_n34), .ZN(u4_sll_482_n35) );
  INV_X4 u4_sll_482_U31 ( .A(u4_sll_482_n33), .ZN(u4_sll_482_n32) );
  INV_X4 u4_sll_482_U30 ( .A(u4_sll_482_n2), .ZN(u4_sll_482_n28) );
  INV_X4 u4_sll_482_U29 ( .A(u4_sll_482_n2), .ZN(u4_sll_482_n24) );
  INV_X4 u4_sll_482_U28 ( .A(u4_sll_482_n2), .ZN(u4_sll_482_n23) );
  INV_X4 u4_sll_482_U27 ( .A(u4_sll_482_n2), .ZN(u4_sll_482_n29) );
  INV_X4 u4_sll_482_U26 ( .A(u4_sll_482_n2), .ZN(u4_sll_482_n25) );
  INV_X4 u4_sll_482_U25 ( .A(u4_sll_482_n12), .ZN(u4_sll_482_n11) );
  INV_X4 u4_sll_482_U24 ( .A(u4_sll_482_temp_int_SH_4_), .ZN(u4_sll_482_n34)
         );
  INV_X4 u4_sll_482_U23 ( .A(u4_sll_482_n1), .ZN(u4_sll_482_n17) );
  INV_X4 u4_sll_482_U22 ( .A(u4_sll_482_n1), .ZN(u4_sll_482_n18) );
  INV_X4 u4_sll_482_U21 ( .A(u4_sll_482_n1), .ZN(u4_sll_482_n15) );
  INV_X4 u4_sll_482_U20 ( .A(u4_sll_482_n33), .ZN(u4_sll_482_n30) );
  INV_X4 u4_sll_482_U19 ( .A(u4_sll_482_n33), .ZN(u4_sll_482_n31) );
  INV_X4 u4_sll_482_U18 ( .A(u4_sll_482_temp_int_SH_3_), .ZN(u4_sll_482_n33)
         );
  AND2_X4 u4_sll_482_U17 ( .A1(u4_sll_482_n19), .A2(u4_sll_482_ML_int_1__113_), 
        .ZN(u4_sll_482_n3) );
  INV_X4 u4_sll_482_U16 ( .A(u4_sll_482_n1), .ZN(u4_sll_482_n20) );
  INV_X4 u4_sll_482_U15 ( .A(u4_sll_482_n1), .ZN(u4_sll_482_n19) );
  INV_X4 u4_sll_482_U14 ( .A(u4_sll_482_n1), .ZN(u4_sll_482_n16) );
  INV_X4 u4_sll_482_U13 ( .A(u4_sll_482_n11), .ZN(u4_sll_482_n6) );
  INV_X4 u4_sll_482_U12 ( .A(u4_sll_482_n2), .ZN(u4_sll_482_n26) );
  INV_X4 u4_sll_482_U11 ( .A(u4_sll_482_n14), .ZN(u4_sll_482_n8) );
  INV_X4 u4_sll_482_U10 ( .A(u4_sll_482_n14), .ZN(u4_sll_482_n12) );
  INV_X4 u4_sll_482_U9 ( .A(u4_sll_482_n10), .ZN(u4_sll_482_n9) );
  INV_X4 u4_sll_482_U8 ( .A(u4_sll_482_temp_int_SH_0_), .ZN(u4_sll_482_n10) );
  INV_X4 u4_sll_482_U7 ( .A(u4_sll_482_n10), .ZN(u4_sll_482_n7) );
  INV_X4 u4_sll_482_U6 ( .A(u4_sll_482_n2), .ZN(u4_sll_482_n27) );
  INV_X4 u4_sll_482_U5 ( .A(u4_sll_482_temp_int_SH_0_), .ZN(u4_sll_482_n14) );
  AND2_X4 u4_sll_482_U4 ( .A1(u4_sll_482_n46), .A2(u4_sll_482_n53), .ZN(
        u4_sll_482_n2) );
  AND2_X4 u4_sll_482_U3 ( .A1(u4_sll_482_n46), .A2(u4_sll_482_n54), .ZN(
        u4_sll_482_n1) );
  MUX2_X2 u4_sll_482_M1_0_1 ( .A(n6344), .B(n6446), .S(u4_sll_482_n13), .Z(
        u4_sll_482_ML_int_1__1_) );
  MUX2_X2 u4_sll_482_M1_0_2 ( .A(n6345), .B(n6344), .S(u4_sll_482_n13), .Z(
        u4_sll_482_ML_int_1__2_) );
  MUX2_X2 u4_sll_482_M1_0_3 ( .A(n6346), .B(n6345), .S(u4_sll_482_n13), .Z(
        u4_sll_482_ML_int_1__3_) );
  MUX2_X2 u4_sll_482_M1_0_4 ( .A(n6347), .B(n6346), .S(u4_sll_482_n9), .Z(
        u4_sll_482_ML_int_1__4_) );
  MUX2_X2 u4_sll_482_M1_0_5 ( .A(n6348), .B(n6347), .S(u4_sll_482_n9), .Z(
        u4_sll_482_ML_int_1__5_) );
  MUX2_X2 u4_sll_482_M1_0_6 ( .A(n6349), .B(n6348), .S(u4_sll_482_n9), .Z(
        u4_sll_482_ML_int_1__6_) );
  MUX2_X2 u4_sll_482_M1_0_7 ( .A(n6350), .B(n6349), .S(u4_sll_482_n9), .Z(
        u4_sll_482_ML_int_1__7_) );
  MUX2_X2 u4_sll_482_M1_0_8 ( .A(n6351), .B(n6350), .S(u4_sll_482_n9), .Z(
        u4_sll_482_ML_int_1__8_) );
  MUX2_X2 u4_sll_482_M1_0_9 ( .A(n6444), .B(n6351), .S(u4_sll_482_n9), .Z(
        u4_sll_482_ML_int_1__9_) );
  MUX2_X2 u4_sll_482_M1_0_10 ( .A(n6443), .B(n6444), .S(u4_sll_482_n9), .Z(
        u4_sll_482_ML_int_1__10_) );
  MUX2_X2 u4_sll_482_M1_0_11 ( .A(n6411), .B(n6443), .S(u4_sll_482_n9), .Z(
        u4_sll_482_ML_int_1__11_) );
  MUX2_X2 u4_sll_482_M1_0_12 ( .A(n6413), .B(n6411), .S(u4_sll_482_n9), .Z(
        u4_sll_482_ML_int_1__12_) );
  MUX2_X2 u4_sll_482_M1_0_13 ( .A(n6414), .B(n6413), .S(u4_sll_482_n9), .Z(
        u4_sll_482_ML_int_1__13_) );
  MUX2_X2 u4_sll_482_M1_0_14 ( .A(n6415), .B(n6414), .S(u4_sll_482_n9), .Z(
        u4_sll_482_ML_int_1__14_) );
  MUX2_X2 u4_sll_482_M1_0_15 ( .A(n6418), .B(n6415), .S(u4_sll_482_n6), .Z(
        u4_sll_482_ML_int_1__15_) );
  MUX2_X2 u4_sll_482_M1_0_16 ( .A(n6416), .B(n6418), .S(u4_sll_482_n13), .Z(
        u4_sll_482_ML_int_1__16_) );
  MUX2_X2 u4_sll_482_M1_0_17 ( .A(n6417), .B(n6416), .S(u4_sll_482_n7), .Z(
        u4_sll_482_ML_int_1__17_) );
  MUX2_X2 u4_sll_482_M1_0_18 ( .A(n6442), .B(n6417), .S(u4_sll_482_n7), .Z(
        u4_sll_482_ML_int_1__18_) );
  MUX2_X2 u4_sll_482_M1_0_19 ( .A(n6419), .B(n6442), .S(u4_sll_482_n7), .Z(
        u4_sll_482_ML_int_1__19_) );
  MUX2_X2 u4_sll_482_M1_0_20 ( .A(n6420), .B(n6419), .S(u4_sll_482_n7), .Z(
        u4_sll_482_ML_int_1__20_) );
  MUX2_X2 u4_sll_482_M1_0_21 ( .A(n6421), .B(n6420), .S(u4_sll_482_n7), .Z(
        u4_sll_482_ML_int_1__21_) );
  MUX2_X2 u4_sll_482_M1_0_22 ( .A(n6422), .B(n6421), .S(u4_sll_482_n7), .Z(
        u4_sll_482_ML_int_1__22_) );
  MUX2_X2 u4_sll_482_M1_0_23 ( .A(n6425), .B(n6422), .S(u4_sll_482_n7), .Z(
        u4_sll_482_ML_int_1__23_) );
  MUX2_X2 u4_sll_482_M1_0_24 ( .A(n6423), .B(n6425), .S(u4_sll_482_n13), .Z(
        u4_sll_482_ML_int_1__24_) );
  MUX2_X2 u4_sll_482_M1_0_25 ( .A(n6424), .B(n6423), .S(u4_sll_482_n7), .Z(
        u4_sll_482_ML_int_1__25_) );
  MUX2_X2 u4_sll_482_M1_0_26 ( .A(n6441), .B(n6424), .S(u4_sll_482_n8), .Z(
        u4_sll_482_ML_int_1__26_) );
  MUX2_X2 u4_sll_482_M1_0_27 ( .A(n6426), .B(n6441), .S(u4_sll_482_n8), .Z(
        u4_sll_482_ML_int_1__27_) );
  MUX2_X2 u4_sll_482_M1_0_28 ( .A(n6427), .B(n6426), .S(u4_sll_482_n8), .Z(
        u4_sll_482_ML_int_1__28_) );
  MUX2_X2 u4_sll_482_M1_0_29 ( .A(n6428), .B(n6427), .S(u4_sll_482_n8), .Z(
        u4_sll_482_ML_int_1__29_) );
  MUX2_X2 u4_sll_482_M1_0_30 ( .A(n6429), .B(n6428), .S(u4_sll_482_n8), .Z(
        u4_sll_482_ML_int_1__30_) );
  MUX2_X2 u4_sll_482_M1_0_31 ( .A(n6432), .B(n6429), .S(u4_sll_482_n8), .Z(
        u4_sll_482_ML_int_1__31_) );
  MUX2_X2 u4_sll_482_M1_0_32 ( .A(n6430), .B(n6432), .S(u4_sll_482_n8), .Z(
        u4_sll_482_ML_int_1__32_) );
  MUX2_X2 u4_sll_482_M1_0_33 ( .A(n6431), .B(n6430), .S(u4_sll_482_n8), .Z(
        u4_sll_482_ML_int_1__33_) );
  MUX2_X2 u4_sll_482_M1_0_34 ( .A(n6440), .B(n6431), .S(u4_sll_482_n8), .Z(
        u4_sll_482_ML_int_1__34_) );
  MUX2_X2 u4_sll_482_M1_0_35 ( .A(n6433), .B(n6440), .S(u4_sll_482_n8), .Z(
        u4_sll_482_ML_int_1__35_) );
  MUX2_X2 u4_sll_482_M1_0_36 ( .A(n6434), .B(n6433), .S(u4_sll_482_n8), .Z(
        u4_sll_482_ML_int_1__36_) );
  MUX2_X2 u4_sll_482_M1_0_37 ( .A(n6435), .B(n6434), .S(u4_sll_482_n13), .Z(
        u4_sll_482_ML_int_1__37_) );
  MUX2_X2 u4_sll_482_M1_0_38 ( .A(n6436), .B(n6435), .S(u4_sll_482_n13), .Z(
        u4_sll_482_ML_int_1__38_) );
  MUX2_X2 u4_sll_482_M1_0_39 ( .A(n6439), .B(n6436), .S(u4_sll_482_n13), .Z(
        u4_sll_482_ML_int_1__39_) );
  MUX2_X2 u4_sll_482_M1_0_40 ( .A(n6437), .B(n6439), .S(u4_sll_482_n13), .Z(
        u4_sll_482_ML_int_1__40_) );
  MUX2_X2 u4_sll_482_M1_0_41 ( .A(n6438), .B(n6437), .S(u4_sll_482_n13), .Z(
        u4_sll_482_ML_int_1__41_) );
  MUX2_X2 u4_sll_482_M1_0_42 ( .A(n6445), .B(n6438), .S(u4_sll_482_n6), .Z(
        u4_sll_482_ML_int_1__42_) );
  MUX2_X2 u4_sll_482_M1_0_43 ( .A(n6405), .B(n6445), .S(u4_sll_482_n6), .Z(
        u4_sll_482_ML_int_1__43_) );
  MUX2_X2 u4_sll_482_M1_0_44 ( .A(n6406), .B(n6405), .S(u4_sll_482_n13), .Z(
        u4_sll_482_ML_int_1__44_) );
  MUX2_X2 u4_sll_482_M1_0_45 ( .A(n6407), .B(n6406), .S(u4_sll_482_n13), .Z(
        u4_sll_482_ML_int_1__45_) );
  MUX2_X2 u4_sll_482_M1_0_46 ( .A(n6408), .B(n6407), .S(u4_sll_482_n6), .Z(
        u4_sll_482_ML_int_1__46_) );
  MUX2_X2 u4_sll_482_M1_0_47 ( .A(n6410), .B(n6408), .S(u4_sll_482_n13), .Z(
        u4_sll_482_ML_int_1__47_) );
  MUX2_X2 u4_sll_482_M1_0_48 ( .A(n6409), .B(n6410), .S(u4_sll_482_n7), .Z(
        u4_sll_482_ML_int_1__48_) );
  MUX2_X2 u4_sll_482_M1_0_49 ( .A(n6367), .B(n6409), .S(u4_sll_482_n7), .Z(
        u4_sll_482_ML_int_1__49_) );
  MUX2_X2 u4_sll_482_M1_0_50 ( .A(fract_denorm[50]), .B(n6367), .S(
        u4_sll_482_n7), .Z(u4_sll_482_ML_int_1__50_) );
  MUX2_X2 u4_sll_482_M1_0_51 ( .A(fract_denorm[51]), .B(fract_denorm[50]), .S(
        u4_sll_482_n7), .Z(u4_sll_482_ML_int_1__51_) );
  MUX2_X2 u4_sll_482_M1_0_52 ( .A(fract_denorm[52]), .B(fract_denorm[51]), .S(
        u4_sll_482_n7), .Z(u4_sll_482_ML_int_1__52_) );
  MUX2_X2 u4_sll_482_M1_0_53 ( .A(fract_denorm[53]), .B(fract_denorm[52]), .S(
        u4_sll_482_n7), .Z(u4_sll_482_ML_int_1__53_) );
  MUX2_X2 u4_sll_482_M1_0_54 ( .A(fract_denorm[54]), .B(fract_denorm[53]), .S(
        u4_sll_482_n7), .Z(u4_sll_482_ML_int_1__54_) );
  MUX2_X2 u4_sll_482_M1_0_55 ( .A(fract_denorm[55]), .B(fract_denorm[54]), .S(
        u4_sll_482_n7), .Z(u4_sll_482_ML_int_1__55_) );
  MUX2_X2 u4_sll_482_M1_0_56 ( .A(fract_denorm[56]), .B(fract_denorm[55]), .S(
        u4_sll_482_n7), .Z(u4_sll_482_ML_int_1__56_) );
  MUX2_X2 u4_sll_482_M1_0_57 ( .A(fract_denorm[57]), .B(fract_denorm[56]), .S(
        u4_sll_482_n7), .Z(u4_sll_482_ML_int_1__57_) );
  MUX2_X2 u4_sll_482_M1_0_58 ( .A(fract_denorm[58]), .B(fract_denorm[57]), .S(
        u4_sll_482_n7), .Z(u4_sll_482_ML_int_1__58_) );
  MUX2_X2 u4_sll_482_M1_0_59 ( .A(fract_denorm[59]), .B(fract_denorm[58]), .S(
        u4_sll_482_n9), .Z(u4_sll_482_ML_int_1__59_) );
  MUX2_X2 u4_sll_482_M1_0_60 ( .A(fract_denorm[60]), .B(fract_denorm[59]), .S(
        u4_sll_482_n12), .Z(u4_sll_482_ML_int_1__60_) );
  MUX2_X2 u4_sll_482_M1_0_61 ( .A(fract_denorm[61]), .B(fract_denorm[60]), .S(
        u4_sll_482_n13), .Z(u4_sll_482_ML_int_1__61_) );
  MUX2_X2 u4_sll_482_M1_0_62 ( .A(fract_denorm[62]), .B(fract_denorm[61]), .S(
        u4_sll_482_n12), .Z(u4_sll_482_ML_int_1__62_) );
  MUX2_X2 u4_sll_482_M1_0_63 ( .A(fract_denorm[63]), .B(fract_denorm[62]), .S(
        u4_sll_482_n12), .Z(u4_sll_482_ML_int_1__63_) );
  MUX2_X2 u4_sll_482_M1_0_64 ( .A(fract_denorm[64]), .B(fract_denorm[63]), .S(
        u4_sll_482_n9), .Z(u4_sll_482_ML_int_1__64_) );
  MUX2_X2 u4_sll_482_M1_0_65 ( .A(fract_denorm[65]), .B(fract_denorm[64]), .S(
        u4_sll_482_n13), .Z(u4_sll_482_ML_int_1__65_) );
  MUX2_X2 u4_sll_482_M1_0_66 ( .A(fract_denorm[66]), .B(fract_denorm[65]), .S(
        u4_sll_482_n8), .Z(u4_sll_482_ML_int_1__66_) );
  MUX2_X2 u4_sll_482_M1_0_67 ( .A(fract_denorm[67]), .B(fract_denorm[66]), .S(
        u4_sll_482_n13), .Z(u4_sll_482_ML_int_1__67_) );
  MUX2_X2 u4_sll_482_M1_0_68 ( .A(fract_denorm[68]), .B(fract_denorm[67]), .S(
        u4_sll_482_n12), .Z(u4_sll_482_ML_int_1__68_) );
  MUX2_X2 u4_sll_482_M1_0_69 ( .A(fract_denorm[69]), .B(fract_denorm[68]), .S(
        u4_sll_482_n12), .Z(u4_sll_482_ML_int_1__69_) );
  MUX2_X2 u4_sll_482_M1_0_70 ( .A(fract_denorm[70]), .B(fract_denorm[69]), .S(
        u4_sll_482_n8), .Z(u4_sll_482_ML_int_1__70_) );
  MUX2_X2 u4_sll_482_M1_0_71 ( .A(fract_denorm[71]), .B(fract_denorm[70]), .S(
        u4_sll_482_n8), .Z(u4_sll_482_ML_int_1__71_) );
  MUX2_X2 u4_sll_482_M1_0_72 ( .A(fract_denorm[72]), .B(fract_denorm[71]), .S(
        u4_sll_482_n8), .Z(u4_sll_482_ML_int_1__72_) );
  MUX2_X2 u4_sll_482_M1_0_73 ( .A(fract_denorm[73]), .B(fract_denorm[72]), .S(
        u4_sll_482_n8), .Z(u4_sll_482_ML_int_1__73_) );
  MUX2_X2 u4_sll_482_M1_0_74 ( .A(fract_denorm[74]), .B(fract_denorm[73]), .S(
        u4_sll_482_n8), .Z(u4_sll_482_ML_int_1__74_) );
  MUX2_X2 u4_sll_482_M1_0_75 ( .A(fract_denorm[75]), .B(fract_denorm[74]), .S(
        u4_sll_482_n8), .Z(u4_sll_482_ML_int_1__75_) );
  MUX2_X2 u4_sll_482_M1_0_76 ( .A(fract_denorm[76]), .B(fract_denorm[75]), .S(
        u4_sll_482_n13), .Z(u4_sll_482_ML_int_1__76_) );
  MUX2_X2 u4_sll_482_M1_0_77 ( .A(fract_denorm[77]), .B(fract_denorm[76]), .S(
        u4_sll_482_n8), .Z(u4_sll_482_ML_int_1__77_) );
  MUX2_X2 u4_sll_482_M1_0_78 ( .A(fract_denorm[78]), .B(fract_denorm[77]), .S(
        u4_sll_482_n13), .Z(u4_sll_482_ML_int_1__78_) );
  MUX2_X2 u4_sll_482_M1_0_79 ( .A(fract_denorm[79]), .B(fract_denorm[78]), .S(
        u4_sll_482_n8), .Z(u4_sll_482_ML_int_1__79_) );
  MUX2_X2 u4_sll_482_M1_0_80 ( .A(fract_denorm[80]), .B(fract_denorm[79]), .S(
        u4_sll_482_n8), .Z(u4_sll_482_ML_int_1__80_) );
  MUX2_X2 u4_sll_482_M1_0_81 ( .A(fract_denorm[81]), .B(fract_denorm[80]), .S(
        u4_sll_482_n13), .Z(u4_sll_482_ML_int_1__81_) );
  MUX2_X2 u4_sll_482_M1_0_82 ( .A(fract_denorm[82]), .B(fract_denorm[81]), .S(
        u4_sll_482_n9), .Z(u4_sll_482_ML_int_1__82_) );
  MUX2_X2 u4_sll_482_M1_0_83 ( .A(fract_denorm[83]), .B(fract_denorm[82]), .S(
        u4_sll_482_n9), .Z(u4_sll_482_ML_int_1__83_) );
  MUX2_X2 u4_sll_482_M1_0_84 ( .A(fract_denorm[84]), .B(fract_denorm[83]), .S(
        u4_sll_482_n12), .Z(u4_sll_482_ML_int_1__84_) );
  MUX2_X2 u4_sll_482_M1_0_85 ( .A(fract_denorm[85]), .B(fract_denorm[84]), .S(
        u4_sll_482_n12), .Z(u4_sll_482_ML_int_1__85_) );
  MUX2_X2 u4_sll_482_M1_0_86 ( .A(fract_denorm[86]), .B(fract_denorm[85]), .S(
        u4_sll_482_n13), .Z(u4_sll_482_ML_int_1__86_) );
  MUX2_X2 u4_sll_482_M1_0_87 ( .A(fract_denorm[87]), .B(fract_denorm[86]), .S(
        u4_sll_482_n13), .Z(u4_sll_482_ML_int_1__87_) );
  MUX2_X2 u4_sll_482_M1_0_88 ( .A(fract_denorm[88]), .B(fract_denorm[87]), .S(
        u4_sll_482_n13), .Z(u4_sll_482_ML_int_1__88_) );
  MUX2_X2 u4_sll_482_M1_0_89 ( .A(fract_denorm[89]), .B(fract_denorm[88]), .S(
        u4_sll_482_n9), .Z(u4_sll_482_ML_int_1__89_) );
  MUX2_X2 u4_sll_482_M1_0_90 ( .A(fract_denorm[90]), .B(fract_denorm[89]), .S(
        u4_sll_482_n12), .Z(u4_sll_482_ML_int_1__90_) );
  MUX2_X2 u4_sll_482_M1_0_91 ( .A(fract_denorm[91]), .B(fract_denorm[90]), .S(
        u4_sll_482_n12), .Z(u4_sll_482_ML_int_1__91_) );
  MUX2_X2 u4_sll_482_M1_0_92 ( .A(fract_denorm[92]), .B(fract_denorm[91]), .S(
        u4_sll_482_n13), .Z(u4_sll_482_ML_int_1__92_) );
  MUX2_X2 u4_sll_482_M1_0_93 ( .A(fract_denorm[93]), .B(fract_denorm[92]), .S(
        u4_sll_482_n13), .Z(u4_sll_482_ML_int_1__93_) );
  MUX2_X2 u4_sll_482_M1_0_94 ( .A(fract_denorm[94]), .B(fract_denorm[93]), .S(
        u4_sll_482_n6), .Z(u4_sll_482_ML_int_1__94_) );
  MUX2_X2 u4_sll_482_M1_0_95 ( .A(fract_denorm[95]), .B(fract_denorm[94]), .S(
        u4_sll_482_n8), .Z(u4_sll_482_ML_int_1__95_) );
  MUX2_X2 u4_sll_482_M1_0_96 ( .A(fract_denorm[96]), .B(fract_denorm[95]), .S(
        u4_sll_482_n8), .Z(u4_sll_482_ML_int_1__96_) );
  MUX2_X2 u4_sll_482_M1_0_97 ( .A(fract_denorm[97]), .B(fract_denorm[96]), .S(
        u4_sll_482_n6), .Z(u4_sll_482_ML_int_1__97_) );
  MUX2_X2 u4_sll_482_M1_0_98 ( .A(fract_denorm[98]), .B(fract_denorm[97]), .S(
        u4_sll_482_n8), .Z(u4_sll_482_ML_int_1__98_) );
  MUX2_X2 u4_sll_482_M1_0_99 ( .A(fract_denorm[99]), .B(fract_denorm[98]), .S(
        u4_sll_482_n6), .Z(u4_sll_482_ML_int_1__99_) );
  MUX2_X2 u4_sll_482_M1_0_100 ( .A(fract_denorm[100]), .B(fract_denorm[99]), 
        .S(u4_sll_482_n13), .Z(u4_sll_482_ML_int_1__100_) );
  MUX2_X2 u4_sll_482_M1_0_101 ( .A(fract_denorm[101]), .B(fract_denorm[100]), 
        .S(u4_sll_482_n13), .Z(u4_sll_482_ML_int_1__101_) );
  MUX2_X2 u4_sll_482_M1_0_102 ( .A(fract_denorm[102]), .B(fract_denorm[101]), 
        .S(u4_sll_482_n8), .Z(u4_sll_482_ML_int_1__102_) );
  MUX2_X2 u4_sll_482_M1_0_103 ( .A(fract_denorm[103]), .B(fract_denorm[102]), 
        .S(u4_sll_482_n6), .Z(u4_sll_482_ML_int_1__103_) );
  MUX2_X2 u4_sll_482_M1_0_104 ( .A(fract_denorm[104]), .B(fract_denorm[103]), 
        .S(u4_sll_482_n6), .Z(u4_sll_482_ML_int_1__104_) );
  MUX2_X2 u4_sll_482_M1_0_105 ( .A(fract_denorm[105]), .B(fract_denorm[104]), 
        .S(u4_sll_482_n6), .Z(u4_sll_482_ML_int_1__105_) );
  MUX2_X2 u4_sll_482_M1_0_106 ( .A(fract_denorm[105]), .B(fract_denorm[105]), 
        .S(u4_sll_482_n6), .Z(u4_sll_482_ML_int_1__106_) );
  MUX2_X2 u4_sll_482_M1_0_107 ( .A(n4652), .B(fract_denorm[105]), .S(
        u4_sll_482_n6), .Z(u4_sll_482_ML_int_1__107_) );
  MUX2_X2 u4_sll_482_M1_0_108 ( .A(n4652), .B(n4652), .S(u4_sll_482_n6), .Z(
        u4_sll_482_ML_int_1__108_) );
  MUX2_X2 u4_sll_482_M1_0_109 ( .A(fract_denorm[105]), .B(n4652), .S(
        u4_sll_482_n6), .Z(u4_sll_482_ML_int_1__109_) );
  MUX2_X2 u4_sll_482_M1_0_110 ( .A(fract_denorm[105]), .B(fract_denorm[105]), 
        .S(u4_sll_482_n6), .Z(u4_sll_482_ML_int_1__110_) );
  MUX2_X2 u4_sll_482_M1_0_111 ( .A(fract_denorm[105]), .B(fract_denorm[105]), 
        .S(u4_sll_482_n6), .Z(u4_sll_482_ML_int_1__111_) );
  MUX2_X2 u4_sll_482_M1_0_112 ( .A(fract_denorm[105]), .B(fract_denorm[105]), 
        .S(u4_sll_482_n6), .Z(u4_sll_482_ML_int_1__112_) );
  MUX2_X2 u4_sll_482_M1_0_113 ( .A(fract_denorm[105]), .B(fract_denorm[105]), 
        .S(u4_sll_482_n6), .Z(u4_sll_482_ML_int_1__113_) );
  MUX2_X2 u4_sll_482_M1_1_2 ( .A(u4_sll_482_ML_int_1__2_), .B(
        u4_sll_482_ML_int_1__0_), .S(u4_sll_482_n15), .Z(
        u4_sll_482_ML_int_2__2_) );
  MUX2_X2 u4_sll_482_M1_1_3 ( .A(u4_sll_482_ML_int_1__3_), .B(
        u4_sll_482_ML_int_1__1_), .S(u4_sll_482_n15), .Z(
        u4_sll_482_ML_int_2__3_) );
  MUX2_X2 u4_sll_482_M1_1_4 ( .A(u4_sll_482_ML_int_1__4_), .B(
        u4_sll_482_ML_int_1__2_), .S(u4_sll_482_n15), .Z(
        u4_sll_482_ML_int_2__4_) );
  MUX2_X2 u4_sll_482_M1_1_5 ( .A(u4_sll_482_ML_int_1__5_), .B(
        u4_sll_482_ML_int_1__3_), .S(u4_sll_482_n15), .Z(
        u4_sll_482_ML_int_2__5_) );
  MUX2_X2 u4_sll_482_M1_1_6 ( .A(u4_sll_482_ML_int_1__6_), .B(
        u4_sll_482_ML_int_1__4_), .S(u4_sll_482_n15), .Z(
        u4_sll_482_ML_int_2__6_) );
  MUX2_X2 u4_sll_482_M1_1_7 ( .A(u4_sll_482_ML_int_1__7_), .B(
        u4_sll_482_ML_int_1__5_), .S(u4_sll_482_n15), .Z(
        u4_sll_482_ML_int_2__7_) );
  MUX2_X2 u4_sll_482_M1_1_8 ( .A(u4_sll_482_ML_int_1__8_), .B(
        u4_sll_482_ML_int_1__6_), .S(u4_sll_482_n15), .Z(
        u4_sll_482_ML_int_2__8_) );
  MUX2_X2 u4_sll_482_M1_1_9 ( .A(u4_sll_482_ML_int_1__9_), .B(
        u4_sll_482_ML_int_1__7_), .S(u4_sll_482_n15), .Z(
        u4_sll_482_ML_int_2__9_) );
  MUX2_X2 u4_sll_482_M1_1_10 ( .A(u4_sll_482_ML_int_1__10_), .B(
        u4_sll_482_ML_int_1__8_), .S(u4_sll_482_n15), .Z(
        u4_sll_482_ML_int_2__10_) );
  MUX2_X2 u4_sll_482_M1_1_11 ( .A(u4_sll_482_ML_int_1__11_), .B(
        u4_sll_482_ML_int_1__9_), .S(u4_sll_482_n15), .Z(
        u4_sll_482_ML_int_2__11_) );
  MUX2_X2 u4_sll_482_M1_1_12 ( .A(u4_sll_482_ML_int_1__12_), .B(
        u4_sll_482_ML_int_1__10_), .S(u4_sll_482_n15), .Z(
        u4_sll_482_ML_int_2__12_) );
  MUX2_X2 u4_sll_482_M1_1_13 ( .A(u4_sll_482_ML_int_1__13_), .B(
        u4_sll_482_ML_int_1__11_), .S(u4_sll_482_n17), .Z(
        u4_sll_482_ML_int_2__13_) );
  MUX2_X2 u4_sll_482_M1_1_14 ( .A(u4_sll_482_ML_int_1__14_), .B(
        u4_sll_482_ML_int_1__12_), .S(u4_sll_482_n17), .Z(
        u4_sll_482_ML_int_2__14_) );
  MUX2_X2 u4_sll_482_M1_1_15 ( .A(u4_sll_482_ML_int_1__15_), .B(
        u4_sll_482_ML_int_1__13_), .S(u4_sll_482_n20), .Z(
        u4_sll_482_ML_int_2__15_) );
  MUX2_X2 u4_sll_482_M1_1_16 ( .A(u4_sll_482_ML_int_1__16_), .B(
        u4_sll_482_ML_int_1__14_), .S(u4_sll_482_n18), .Z(
        u4_sll_482_ML_int_2__16_) );
  MUX2_X2 u4_sll_482_M1_1_17 ( .A(u4_sll_482_ML_int_1__17_), .B(
        u4_sll_482_ML_int_1__15_), .S(u4_sll_482_n20), .Z(
        u4_sll_482_ML_int_2__17_) );
  MUX2_X2 u4_sll_482_M1_1_18 ( .A(u4_sll_482_ML_int_1__18_), .B(
        u4_sll_482_ML_int_1__16_), .S(u4_sll_482_n16), .Z(
        u4_sll_482_ML_int_2__18_) );
  MUX2_X2 u4_sll_482_M1_1_19 ( .A(u4_sll_482_ML_int_1__19_), .B(
        u4_sll_482_ML_int_1__17_), .S(u4_sll_482_n18), .Z(
        u4_sll_482_ML_int_2__19_) );
  MUX2_X2 u4_sll_482_M1_1_20 ( .A(u4_sll_482_ML_int_1__20_), .B(
        u4_sll_482_ML_int_1__18_), .S(u4_sll_482_n16), .Z(
        u4_sll_482_ML_int_2__20_) );
  MUX2_X2 u4_sll_482_M1_1_21 ( .A(u4_sll_482_ML_int_1__21_), .B(
        u4_sll_482_ML_int_1__19_), .S(u4_sll_482_n19), .Z(
        u4_sll_482_ML_int_2__21_) );
  MUX2_X2 u4_sll_482_M1_1_22 ( .A(u4_sll_482_ML_int_1__22_), .B(
        u4_sll_482_ML_int_1__20_), .S(u4_sll_482_n15), .Z(
        u4_sll_482_ML_int_2__22_) );
  MUX2_X2 u4_sll_482_M1_1_23 ( .A(u4_sll_482_ML_int_1__23_), .B(
        u4_sll_482_ML_int_1__21_), .S(u4_sll_482_n15), .Z(
        u4_sll_482_ML_int_2__23_) );
  MUX2_X2 u4_sll_482_M1_1_24 ( .A(u4_sll_482_ML_int_1__24_), .B(
        u4_sll_482_ML_int_1__22_), .S(u4_sll_482_n16), .Z(
        u4_sll_482_ML_int_2__24_) );
  MUX2_X2 u4_sll_482_M1_1_25 ( .A(u4_sll_482_ML_int_1__25_), .B(
        u4_sll_482_ML_int_1__23_), .S(u4_sll_482_n16), .Z(
        u4_sll_482_ML_int_2__25_) );
  MUX2_X2 u4_sll_482_M1_1_26 ( .A(u4_sll_482_ML_int_1__26_), .B(
        u4_sll_482_ML_int_1__24_), .S(u4_sll_482_n16), .Z(
        u4_sll_482_ML_int_2__26_) );
  MUX2_X2 u4_sll_482_M1_1_27 ( .A(u4_sll_482_ML_int_1__27_), .B(
        u4_sll_482_ML_int_1__25_), .S(u4_sll_482_n16), .Z(
        u4_sll_482_ML_int_2__27_) );
  MUX2_X2 u4_sll_482_M1_1_28 ( .A(u4_sll_482_ML_int_1__28_), .B(
        u4_sll_482_ML_int_1__26_), .S(u4_sll_482_n16), .Z(
        u4_sll_482_ML_int_2__28_) );
  MUX2_X2 u4_sll_482_M1_1_29 ( .A(u4_sll_482_ML_int_1__29_), .B(
        u4_sll_482_ML_int_1__27_), .S(u4_sll_482_n16), .Z(
        u4_sll_482_ML_int_2__29_) );
  MUX2_X2 u4_sll_482_M1_1_30 ( .A(u4_sll_482_ML_int_1__30_), .B(
        u4_sll_482_ML_int_1__28_), .S(u4_sll_482_n16), .Z(
        u4_sll_482_ML_int_2__30_) );
  MUX2_X2 u4_sll_482_M1_1_31 ( .A(u4_sll_482_ML_int_1__31_), .B(
        u4_sll_482_ML_int_1__29_), .S(u4_sll_482_n16), .Z(
        u4_sll_482_ML_int_2__31_) );
  MUX2_X2 u4_sll_482_M1_1_32 ( .A(u4_sll_482_ML_int_1__32_), .B(
        u4_sll_482_ML_int_1__30_), .S(u4_sll_482_n16), .Z(
        u4_sll_482_ML_int_2__32_) );
  MUX2_X2 u4_sll_482_M1_1_33 ( .A(u4_sll_482_ML_int_1__33_), .B(
        u4_sll_482_ML_int_1__31_), .S(u4_sll_482_n16), .Z(
        u4_sll_482_ML_int_2__33_) );
  MUX2_X2 u4_sll_482_M1_1_34 ( .A(u4_sll_482_ML_int_1__34_), .B(
        u4_sll_482_ML_int_1__32_), .S(u4_sll_482_n16), .Z(
        u4_sll_482_ML_int_2__34_) );
  MUX2_X2 u4_sll_482_M1_1_35 ( .A(u4_sll_482_ML_int_1__35_), .B(
        u4_sll_482_ML_int_1__33_), .S(u4_sll_482_n17), .Z(
        u4_sll_482_ML_int_2__35_) );
  MUX2_X2 u4_sll_482_M1_1_36 ( .A(u4_sll_482_ML_int_1__36_), .B(
        u4_sll_482_ML_int_1__34_), .S(u4_sll_482_n17), .Z(
        u4_sll_482_ML_int_2__36_) );
  MUX2_X2 u4_sll_482_M1_1_37 ( .A(u4_sll_482_ML_int_1__37_), .B(
        u4_sll_482_ML_int_1__35_), .S(u4_sll_482_n17), .Z(
        u4_sll_482_ML_int_2__37_) );
  MUX2_X2 u4_sll_482_M1_1_38 ( .A(u4_sll_482_ML_int_1__38_), .B(
        u4_sll_482_ML_int_1__36_), .S(u4_sll_482_n17), .Z(
        u4_sll_482_ML_int_2__38_) );
  MUX2_X2 u4_sll_482_M1_1_39 ( .A(u4_sll_482_ML_int_1__39_), .B(
        u4_sll_482_ML_int_1__37_), .S(u4_sll_482_n17), .Z(
        u4_sll_482_ML_int_2__39_) );
  MUX2_X2 u4_sll_482_M1_1_40 ( .A(u4_sll_482_ML_int_1__40_), .B(
        u4_sll_482_ML_int_1__38_), .S(u4_sll_482_n17), .Z(
        u4_sll_482_ML_int_2__40_) );
  MUX2_X2 u4_sll_482_M1_1_41 ( .A(u4_sll_482_ML_int_1__41_), .B(
        u4_sll_482_ML_int_1__39_), .S(u4_sll_482_n17), .Z(
        u4_sll_482_ML_int_2__41_) );
  MUX2_X2 u4_sll_482_M1_1_42 ( .A(u4_sll_482_ML_int_1__42_), .B(
        u4_sll_482_ML_int_1__40_), .S(u4_sll_482_n17), .Z(
        u4_sll_482_ML_int_2__42_) );
  MUX2_X2 u4_sll_482_M1_1_43 ( .A(u4_sll_482_ML_int_1__43_), .B(
        u4_sll_482_ML_int_1__41_), .S(u4_sll_482_n17), .Z(
        u4_sll_482_ML_int_2__43_) );
  MUX2_X2 u4_sll_482_M1_1_44 ( .A(u4_sll_482_ML_int_1__44_), .B(
        u4_sll_482_ML_int_1__42_), .S(u4_sll_482_n17), .Z(
        u4_sll_482_ML_int_2__44_) );
  MUX2_X2 u4_sll_482_M1_1_45 ( .A(u4_sll_482_ML_int_1__45_), .B(
        u4_sll_482_ML_int_1__43_), .S(u4_sll_482_n17), .Z(
        u4_sll_482_ML_int_2__45_) );
  MUX2_X2 u4_sll_482_M1_1_46 ( .A(u4_sll_482_ML_int_1__46_), .B(
        u4_sll_482_ML_int_1__44_), .S(u4_sll_482_n20), .Z(
        u4_sll_482_ML_int_2__46_) );
  MUX2_X2 u4_sll_482_M1_1_47 ( .A(u4_sll_482_ML_int_1__47_), .B(
        u4_sll_482_ML_int_1__45_), .S(u4_sll_482_n20), .Z(
        u4_sll_482_ML_int_2__47_) );
  MUX2_X2 u4_sll_482_M1_1_48 ( .A(u4_sll_482_ML_int_1__48_), .B(
        u4_sll_482_ML_int_1__46_), .S(u4_sll_482_n20), .Z(
        u4_sll_482_ML_int_2__48_) );
  MUX2_X2 u4_sll_482_M1_1_49 ( .A(u4_sll_482_ML_int_1__49_), .B(
        u4_sll_482_ML_int_1__47_), .S(u4_sll_482_n20), .Z(
        u4_sll_482_ML_int_2__49_) );
  MUX2_X2 u4_sll_482_M1_1_50 ( .A(u4_sll_482_ML_int_1__50_), .B(
        u4_sll_482_ML_int_1__48_), .S(u4_sll_482_n20), .Z(
        u4_sll_482_ML_int_2__50_) );
  MUX2_X2 u4_sll_482_M1_1_51 ( .A(u4_sll_482_ML_int_1__51_), .B(
        u4_sll_482_ML_int_1__49_), .S(u4_sll_482_n20), .Z(
        u4_sll_482_ML_int_2__51_) );
  MUX2_X2 u4_sll_482_M1_1_52 ( .A(u4_sll_482_ML_int_1__52_), .B(
        u4_sll_482_ML_int_1__50_), .S(u4_sll_482_n20), .Z(
        u4_sll_482_ML_int_2__52_) );
  MUX2_X2 u4_sll_482_M1_1_53 ( .A(u4_sll_482_ML_int_1__53_), .B(
        u4_sll_482_ML_int_1__51_), .S(u4_sll_482_n20), .Z(
        u4_sll_482_ML_int_2__53_) );
  MUX2_X2 u4_sll_482_M1_1_54 ( .A(u4_sll_482_ML_int_1__54_), .B(
        u4_sll_482_ML_int_1__52_), .S(u4_sll_482_n16), .Z(
        u4_sll_482_ML_int_2__54_) );
  MUX2_X2 u4_sll_482_M1_1_55 ( .A(u4_sll_482_ML_int_1__55_), .B(
        u4_sll_482_ML_int_1__53_), .S(u4_sll_482_n19), .Z(
        u4_sll_482_ML_int_2__55_) );
  MUX2_X2 u4_sll_482_M1_1_56 ( .A(u4_sll_482_ML_int_1__56_), .B(
        u4_sll_482_ML_int_1__54_), .S(u4_sll_482_n20), .Z(
        u4_sll_482_ML_int_2__56_) );
  MUX2_X2 u4_sll_482_M1_1_57 ( .A(u4_sll_482_ML_int_1__57_), .B(
        u4_sll_482_ML_int_1__55_), .S(u4_sll_482_n18), .Z(
        u4_sll_482_ML_int_2__57_) );
  MUX2_X2 u4_sll_482_M1_1_58 ( .A(u4_sll_482_ML_int_1__58_), .B(
        u4_sll_482_ML_int_1__56_), .S(u4_sll_482_n18), .Z(
        u4_sll_482_ML_int_2__58_) );
  MUX2_X2 u4_sll_482_M1_1_59 ( .A(u4_sll_482_ML_int_1__59_), .B(
        u4_sll_482_ML_int_1__57_), .S(u4_sll_482_n18), .Z(
        u4_sll_482_ML_int_2__59_) );
  MUX2_X2 u4_sll_482_M1_1_60 ( .A(u4_sll_482_ML_int_1__60_), .B(
        u4_sll_482_ML_int_1__58_), .S(u4_sll_482_n18), .Z(
        u4_sll_482_ML_int_2__60_) );
  MUX2_X2 u4_sll_482_M1_1_61 ( .A(u4_sll_482_ML_int_1__61_), .B(
        u4_sll_482_ML_int_1__59_), .S(u4_sll_482_n18), .Z(
        u4_sll_482_ML_int_2__61_) );
  MUX2_X2 u4_sll_482_M1_1_62 ( .A(u4_sll_482_ML_int_1__62_), .B(
        u4_sll_482_ML_int_1__60_), .S(u4_sll_482_n18), .Z(
        u4_sll_482_ML_int_2__62_) );
  MUX2_X2 u4_sll_482_M1_1_63 ( .A(u4_sll_482_ML_int_1__63_), .B(
        u4_sll_482_ML_int_1__61_), .S(u4_sll_482_n18), .Z(
        u4_sll_482_ML_int_2__63_) );
  MUX2_X2 u4_sll_482_M1_1_64 ( .A(u4_sll_482_ML_int_1__64_), .B(
        u4_sll_482_ML_int_1__62_), .S(u4_sll_482_n18), .Z(
        u4_sll_482_ML_int_2__64_) );
  MUX2_X2 u4_sll_482_M1_1_65 ( .A(u4_sll_482_ML_int_1__65_), .B(
        u4_sll_482_ML_int_1__63_), .S(u4_sll_482_n18), .Z(
        u4_sll_482_ML_int_2__65_) );
  MUX2_X2 u4_sll_482_M1_1_66 ( .A(u4_sll_482_ML_int_1__66_), .B(
        u4_sll_482_ML_int_1__64_), .S(u4_sll_482_n18), .Z(
        u4_sll_482_ML_int_2__66_) );
  MUX2_X2 u4_sll_482_M1_1_67 ( .A(u4_sll_482_ML_int_1__67_), .B(
        u4_sll_482_ML_int_1__65_), .S(u4_sll_482_n18), .Z(
        u4_sll_482_ML_int_2__67_) );
  MUX2_X2 u4_sll_482_M1_1_68 ( .A(u4_sll_482_ML_int_1__68_), .B(
        u4_sll_482_ML_int_1__66_), .S(u4_sll_482_n19), .Z(
        u4_sll_482_ML_int_2__68_) );
  MUX2_X2 u4_sll_482_M1_1_69 ( .A(u4_sll_482_ML_int_1__69_), .B(
        u4_sll_482_ML_int_1__67_), .S(u4_sll_482_n19), .Z(
        u4_sll_482_ML_int_2__69_) );
  MUX2_X2 u4_sll_482_M1_1_70 ( .A(u4_sll_482_ML_int_1__70_), .B(
        u4_sll_482_ML_int_1__68_), .S(u4_sll_482_n19), .Z(
        u4_sll_482_ML_int_2__70_) );
  MUX2_X2 u4_sll_482_M1_1_71 ( .A(u4_sll_482_ML_int_1__71_), .B(
        u4_sll_482_ML_int_1__69_), .S(u4_sll_482_n19), .Z(
        u4_sll_482_ML_int_2__71_) );
  MUX2_X2 u4_sll_482_M1_1_72 ( .A(u4_sll_482_ML_int_1__72_), .B(
        u4_sll_482_ML_int_1__70_), .S(u4_sll_482_n19), .Z(
        u4_sll_482_ML_int_2__72_) );
  MUX2_X2 u4_sll_482_M1_1_73 ( .A(u4_sll_482_ML_int_1__73_), .B(
        u4_sll_482_ML_int_1__71_), .S(u4_sll_482_n19), .Z(
        u4_sll_482_ML_int_2__73_) );
  MUX2_X2 u4_sll_482_M1_1_74 ( .A(u4_sll_482_ML_int_1__74_), .B(
        u4_sll_482_ML_int_1__72_), .S(u4_sll_482_n19), .Z(
        u4_sll_482_ML_int_2__74_) );
  MUX2_X2 u4_sll_482_M1_1_75 ( .A(u4_sll_482_ML_int_1__75_), .B(
        u4_sll_482_ML_int_1__73_), .S(u4_sll_482_n19), .Z(
        u4_sll_482_ML_int_2__75_) );
  MUX2_X2 u4_sll_482_M1_1_76 ( .A(u4_sll_482_ML_int_1__76_), .B(
        u4_sll_482_ML_int_1__74_), .S(u4_sll_482_n19), .Z(
        u4_sll_482_ML_int_2__76_) );
  MUX2_X2 u4_sll_482_M1_1_77 ( .A(u4_sll_482_ML_int_1__77_), .B(
        u4_sll_482_ML_int_1__75_), .S(u4_sll_482_n19), .Z(
        u4_sll_482_ML_int_2__77_) );
  MUX2_X2 u4_sll_482_M1_1_78 ( .A(u4_sll_482_ML_int_1__78_), .B(
        u4_sll_482_ML_int_1__76_), .S(u4_sll_482_n19), .Z(
        u4_sll_482_ML_int_2__78_) );
  MUX2_X2 u4_sll_482_M1_1_79 ( .A(u4_sll_482_ML_int_1__79_), .B(
        u4_sll_482_ML_int_1__77_), .S(u4_sll_482_n20), .Z(
        u4_sll_482_ML_int_2__79_) );
  MUX2_X2 u4_sll_482_M1_1_80 ( .A(u4_sll_482_ML_int_1__80_), .B(
        u4_sll_482_ML_int_1__78_), .S(u4_sll_482_n20), .Z(
        u4_sll_482_ML_int_2__80_) );
  MUX2_X2 u4_sll_482_M1_1_81 ( .A(u4_sll_482_ML_int_1__81_), .B(
        u4_sll_482_ML_int_1__79_), .S(u4_sll_482_n20), .Z(
        u4_sll_482_ML_int_2__81_) );
  MUX2_X2 u4_sll_482_M1_1_82 ( .A(u4_sll_482_ML_int_1__82_), .B(
        u4_sll_482_ML_int_1__80_), .S(u4_sll_482_n20), .Z(
        u4_sll_482_ML_int_2__82_) );
  MUX2_X2 u4_sll_482_M1_1_83 ( .A(u4_sll_482_ML_int_1__83_), .B(
        u4_sll_482_ML_int_1__81_), .S(u4_sll_482_n20), .Z(
        u4_sll_482_ML_int_2__83_) );
  MUX2_X2 u4_sll_482_M1_1_84 ( .A(u4_sll_482_ML_int_1__84_), .B(
        u4_sll_482_ML_int_1__82_), .S(u4_sll_482_n20), .Z(
        u4_sll_482_ML_int_2__84_) );
  MUX2_X2 u4_sll_482_M1_1_85 ( .A(u4_sll_482_ML_int_1__85_), .B(
        u4_sll_482_ML_int_1__83_), .S(u4_sll_482_n20), .Z(
        u4_sll_482_ML_int_2__85_) );
  MUX2_X2 u4_sll_482_M1_1_86 ( .A(u4_sll_482_ML_int_1__86_), .B(
        u4_sll_482_ML_int_1__84_), .S(u4_sll_482_n20), .Z(
        u4_sll_482_ML_int_2__86_) );
  MUX2_X2 u4_sll_482_M1_1_87 ( .A(u4_sll_482_ML_int_1__87_), .B(
        u4_sll_482_ML_int_1__85_), .S(u4_sll_482_n20), .Z(
        u4_sll_482_ML_int_2__87_) );
  MUX2_X2 u4_sll_482_M1_1_88 ( .A(u4_sll_482_ML_int_1__88_), .B(
        u4_sll_482_ML_int_1__86_), .S(u4_sll_482_n20), .Z(
        u4_sll_482_ML_int_2__88_) );
  MUX2_X2 u4_sll_482_M1_1_89 ( .A(u4_sll_482_ML_int_1__89_), .B(
        u4_sll_482_ML_int_1__87_), .S(u4_sll_482_n20), .Z(
        u4_sll_482_ML_int_2__89_) );
  MUX2_X2 u4_sll_482_M1_1_90 ( .A(u4_sll_482_ML_int_1__90_), .B(
        u4_sll_482_ML_int_1__88_), .S(u4_sll_482_n21), .Z(
        u4_sll_482_ML_int_2__90_) );
  MUX2_X2 u4_sll_482_M1_1_91 ( .A(u4_sll_482_ML_int_1__91_), .B(
        u4_sll_482_ML_int_1__89_), .S(u4_sll_482_n21), .Z(
        u4_sll_482_ML_int_2__91_) );
  MUX2_X2 u4_sll_482_M1_1_92 ( .A(u4_sll_482_ML_int_1__92_), .B(
        u4_sll_482_ML_int_1__90_), .S(u4_sll_482_n21), .Z(
        u4_sll_482_ML_int_2__92_) );
  MUX2_X2 u4_sll_482_M1_1_93 ( .A(u4_sll_482_ML_int_1__93_), .B(
        u4_sll_482_ML_int_1__91_), .S(u4_sll_482_n21), .Z(
        u4_sll_482_ML_int_2__93_) );
  MUX2_X2 u4_sll_482_M1_1_94 ( .A(u4_sll_482_ML_int_1__94_), .B(
        u4_sll_482_ML_int_1__92_), .S(u4_sll_482_n21), .Z(
        u4_sll_482_ML_int_2__94_) );
  MUX2_X2 u4_sll_482_M1_1_95 ( .A(u4_sll_482_ML_int_1__95_), .B(
        u4_sll_482_ML_int_1__93_), .S(u4_sll_482_n21), .Z(
        u4_sll_482_ML_int_2__95_) );
  MUX2_X2 u4_sll_482_M1_1_96 ( .A(u4_sll_482_ML_int_1__96_), .B(
        u4_sll_482_ML_int_1__94_), .S(u4_sll_482_n21), .Z(
        u4_sll_482_ML_int_2__96_) );
  MUX2_X2 u4_sll_482_M1_1_97 ( .A(u4_sll_482_ML_int_1__97_), .B(
        u4_sll_482_ML_int_1__95_), .S(u4_sll_482_n21), .Z(
        u4_sll_482_ML_int_2__97_) );
  MUX2_X2 u4_sll_482_M1_1_98 ( .A(u4_sll_482_ML_int_1__98_), .B(
        u4_sll_482_ML_int_1__96_), .S(u4_sll_482_n21), .Z(
        u4_sll_482_ML_int_2__98_) );
  MUX2_X2 u4_sll_482_M1_1_99 ( .A(u4_sll_482_ML_int_1__99_), .B(
        u4_sll_482_ML_int_1__97_), .S(u4_sll_482_n21), .Z(
        u4_sll_482_ML_int_2__99_) );
  MUX2_X2 u4_sll_482_M1_1_100 ( .A(u4_sll_482_ML_int_1__100_), .B(
        u4_sll_482_ML_int_1__98_), .S(u4_sll_482_n21), .Z(
        u4_sll_482_ML_int_2__100_) );
  MUX2_X2 u4_sll_482_M1_1_101 ( .A(u4_sll_482_ML_int_1__101_), .B(
        u4_sll_482_ML_int_1__99_), .S(u4_sll_482_n22), .Z(
        u4_sll_482_ML_int_2__101_) );
  MUX2_X2 u4_sll_482_M1_1_102 ( .A(u4_sll_482_ML_int_1__102_), .B(
        u4_sll_482_ML_int_1__100_), .S(u4_sll_482_n22), .Z(
        u4_sll_482_ML_int_2__102_) );
  MUX2_X2 u4_sll_482_M1_1_103 ( .A(u4_sll_482_ML_int_1__103_), .B(
        u4_sll_482_ML_int_1__101_), .S(u4_sll_482_n22), .Z(
        u4_sll_482_ML_int_2__103_) );
  MUX2_X2 u4_sll_482_M1_1_104 ( .A(u4_sll_482_ML_int_1__104_), .B(
        u4_sll_482_ML_int_1__102_), .S(u4_sll_482_n22), .Z(
        u4_sll_482_ML_int_2__104_) );
  MUX2_X2 u4_sll_482_M1_1_105 ( .A(u4_sll_482_ML_int_1__105_), .B(
        u4_sll_482_ML_int_1__103_), .S(u4_sll_482_n22), .Z(
        u4_sll_482_ML_int_2__105_) );
  MUX2_X2 u4_sll_482_M1_1_106 ( .A(u4_sll_482_ML_int_1__106_), .B(
        u4_sll_482_ML_int_1__104_), .S(u4_sll_482_n22), .Z(
        u4_sll_482_ML_int_2__106_) );
  MUX2_X2 u4_sll_482_M1_1_107 ( .A(u4_sll_482_ML_int_1__107_), .B(
        u4_sll_482_ML_int_1__105_), .S(u4_sll_482_n22), .Z(
        u4_sll_482_ML_int_2__107_) );
  MUX2_X2 u4_sll_482_M1_1_108 ( .A(u4_sll_482_ML_int_1__108_), .B(
        u4_sll_482_ML_int_1__106_), .S(u4_sll_482_n22), .Z(
        u4_sll_482_ML_int_2__108_) );
  MUX2_X2 u4_sll_482_M1_1_109 ( .A(u4_sll_482_ML_int_1__109_), .B(
        u4_sll_482_ML_int_1__107_), .S(u4_sll_482_n22), .Z(
        u4_sll_482_ML_int_2__109_) );
  MUX2_X2 u4_sll_482_M1_1_110 ( .A(u4_sll_482_ML_int_1__110_), .B(
        u4_sll_482_ML_int_1__108_), .S(u4_sll_482_n22), .Z(
        u4_sll_482_ML_int_2__110_) );
  MUX2_X2 u4_sll_482_M1_1_111 ( .A(u4_sll_482_ML_int_1__111_), .B(
        u4_sll_482_ML_int_1__109_), .S(u4_sll_482_n22), .Z(
        u4_sll_482_ML_int_2__111_) );
  MUX2_X2 u4_sll_482_M1_1_112 ( .A(u4_sll_482_ML_int_1__112_), .B(
        u4_sll_482_ML_int_1__110_), .S(u4_sll_482_n19), .Z(
        u4_sll_482_ML_int_2__112_) );
  MUX2_X2 u4_sll_482_M1_1_113 ( .A(u4_sll_482_ML_int_1__113_), .B(
        u4_sll_482_ML_int_1__111_), .S(u4_sll_482_n21), .Z(
        u4_sll_482_ML_int_2__113_) );
  MUX2_X2 u4_sll_482_M1_1_114 ( .A(u4_sll_482_MR_int_1__113_), .B(
        u4_sll_482_ML_int_1__112_), .S(u4_sll_482_n22), .Z(
        u4_sll_482_ML_int_2__114_) );
  MUX2_X2 u4_sll_482_M1_2_4 ( .A(u4_sll_482_ML_int_2__4_), .B(u4_sll_482_n37), 
        .S(u4_sll_482_n23), .Z(u4_sll_482_ML_int_3__4_) );
  MUX2_X2 u4_sll_482_M1_2_5 ( .A(u4_sll_482_ML_int_2__5_), .B(u4_sll_482_n39), 
        .S(u4_sll_482_n23), .Z(u4_sll_482_ML_int_3__5_) );
  MUX2_X2 u4_sll_482_M1_2_6 ( .A(u4_sll_482_ML_int_2__6_), .B(
        u4_sll_482_ML_int_2__2_), .S(u4_sll_482_n23), .Z(
        u4_sll_482_ML_int_3__6_) );
  MUX2_X2 u4_sll_482_M1_2_7 ( .A(u4_sll_482_ML_int_2__7_), .B(
        u4_sll_482_ML_int_2__3_), .S(u4_sll_482_n23), .Z(
        u4_sll_482_ML_int_3__7_) );
  MUX2_X2 u4_sll_482_M1_2_8 ( .A(u4_sll_482_ML_int_2__8_), .B(
        u4_sll_482_ML_int_2__4_), .S(u4_sll_482_n23), .Z(
        u4_sll_482_ML_int_3__8_) );
  MUX2_X2 u4_sll_482_M1_2_9 ( .A(u4_sll_482_ML_int_2__9_), .B(
        u4_sll_482_ML_int_2__5_), .S(u4_sll_482_n23), .Z(
        u4_sll_482_ML_int_3__9_) );
  MUX2_X2 u4_sll_482_M1_2_10 ( .A(u4_sll_482_ML_int_2__10_), .B(
        u4_sll_482_ML_int_2__6_), .S(u4_sll_482_n23), .Z(
        u4_sll_482_ML_int_3__10_) );
  MUX2_X2 u4_sll_482_M1_2_11 ( .A(u4_sll_482_ML_int_2__11_), .B(
        u4_sll_482_ML_int_2__7_), .S(u4_sll_482_n23), .Z(
        u4_sll_482_ML_int_3__11_) );
  MUX2_X2 u4_sll_482_M1_2_12 ( .A(u4_sll_482_ML_int_2__12_), .B(
        u4_sll_482_ML_int_2__8_), .S(u4_sll_482_n23), .Z(
        u4_sll_482_ML_int_3__12_) );
  MUX2_X2 u4_sll_482_M1_2_13 ( .A(u4_sll_482_ML_int_2__13_), .B(
        u4_sll_482_ML_int_2__9_), .S(u4_sll_482_n23), .Z(
        u4_sll_482_ML_int_3__13_) );
  MUX2_X2 u4_sll_482_M1_2_14 ( .A(u4_sll_482_ML_int_2__14_), .B(
        u4_sll_482_ML_int_2__10_), .S(u4_sll_482_n23), .Z(
        u4_sll_482_ML_int_3__14_) );
  MUX2_X2 u4_sll_482_M1_2_15 ( .A(u4_sll_482_ML_int_2__15_), .B(
        u4_sll_482_ML_int_2__11_), .S(u4_sll_482_n24), .Z(
        u4_sll_482_ML_int_3__15_) );
  MUX2_X2 u4_sll_482_M1_2_16 ( .A(u4_sll_482_ML_int_2__16_), .B(
        u4_sll_482_ML_int_2__12_), .S(u4_sll_482_n24), .Z(
        u4_sll_482_ML_int_3__16_) );
  MUX2_X2 u4_sll_482_M1_2_17 ( .A(u4_sll_482_ML_int_2__17_), .B(
        u4_sll_482_ML_int_2__13_), .S(u4_sll_482_n24), .Z(
        u4_sll_482_ML_int_3__17_) );
  MUX2_X2 u4_sll_482_M1_2_18 ( .A(u4_sll_482_ML_int_2__18_), .B(
        u4_sll_482_ML_int_2__14_), .S(u4_sll_482_n24), .Z(
        u4_sll_482_ML_int_3__18_) );
  MUX2_X2 u4_sll_482_M1_2_19 ( .A(u4_sll_482_ML_int_2__19_), .B(
        u4_sll_482_ML_int_2__15_), .S(u4_sll_482_n24), .Z(
        u4_sll_482_ML_int_3__19_) );
  MUX2_X2 u4_sll_482_M1_2_20 ( .A(u4_sll_482_ML_int_2__20_), .B(
        u4_sll_482_ML_int_2__16_), .S(u4_sll_482_n24), .Z(
        u4_sll_482_ML_int_3__20_) );
  MUX2_X2 u4_sll_482_M1_2_21 ( .A(u4_sll_482_ML_int_2__21_), .B(
        u4_sll_482_ML_int_2__17_), .S(u4_sll_482_n24), .Z(
        u4_sll_482_ML_int_3__21_) );
  MUX2_X2 u4_sll_482_M1_2_22 ( .A(u4_sll_482_ML_int_2__22_), .B(
        u4_sll_482_ML_int_2__18_), .S(u4_sll_482_n24), .Z(
        u4_sll_482_ML_int_3__22_) );
  MUX2_X2 u4_sll_482_M1_2_23 ( .A(u4_sll_482_ML_int_2__23_), .B(
        u4_sll_482_ML_int_2__19_), .S(u4_sll_482_n24), .Z(
        u4_sll_482_ML_int_3__23_) );
  MUX2_X2 u4_sll_482_M1_2_24 ( .A(u4_sll_482_ML_int_2__24_), .B(
        u4_sll_482_ML_int_2__20_), .S(u4_sll_482_n24), .Z(
        u4_sll_482_ML_int_3__24_) );
  MUX2_X2 u4_sll_482_M1_2_25 ( .A(u4_sll_482_ML_int_2__25_), .B(
        u4_sll_482_ML_int_2__21_), .S(u4_sll_482_n24), .Z(
        u4_sll_482_ML_int_3__25_) );
  MUX2_X2 u4_sll_482_M1_2_26 ( .A(u4_sll_482_ML_int_2__26_), .B(
        u4_sll_482_ML_int_2__22_), .S(u4_sll_482_n23), .Z(
        u4_sll_482_ML_int_3__26_) );
  MUX2_X2 u4_sll_482_M1_2_27 ( .A(u4_sll_482_ML_int_2__27_), .B(
        u4_sll_482_ML_int_2__23_), .S(u4_sll_482_n24), .Z(
        u4_sll_482_ML_int_3__27_) );
  MUX2_X2 u4_sll_482_M1_2_28 ( .A(u4_sll_482_ML_int_2__28_), .B(
        u4_sll_482_ML_int_2__24_), .S(u4_sll_482_n29), .Z(
        u4_sll_482_ML_int_3__28_) );
  MUX2_X2 u4_sll_482_M1_2_29 ( .A(u4_sll_482_ML_int_2__29_), .B(
        u4_sll_482_ML_int_2__25_), .S(u4_sll_482_n29), .Z(
        u4_sll_482_ML_int_3__29_) );
  MUX2_X2 u4_sll_482_M1_2_30 ( .A(u4_sll_482_ML_int_2__30_), .B(
        u4_sll_482_ML_int_2__26_), .S(u4_sll_482_n29), .Z(
        u4_sll_482_ML_int_3__30_) );
  MUX2_X2 u4_sll_482_M1_2_31 ( .A(u4_sll_482_ML_int_2__31_), .B(
        u4_sll_482_ML_int_2__27_), .S(u4_sll_482_n29), .Z(
        u4_sll_482_ML_int_3__31_) );
  MUX2_X2 u4_sll_482_M1_2_32 ( .A(u4_sll_482_ML_int_2__32_), .B(
        u4_sll_482_ML_int_2__28_), .S(u4_sll_482_n29), .Z(
        u4_sll_482_ML_int_3__32_) );
  MUX2_X2 u4_sll_482_M1_2_33 ( .A(u4_sll_482_ML_int_2__33_), .B(
        u4_sll_482_ML_int_2__29_), .S(u4_sll_482_n29), .Z(
        u4_sll_482_ML_int_3__33_) );
  MUX2_X2 u4_sll_482_M1_2_34 ( .A(u4_sll_482_ML_int_2__34_), .B(
        u4_sll_482_ML_int_2__30_), .S(u4_sll_482_n25), .Z(
        u4_sll_482_ML_int_3__34_) );
  MUX2_X2 u4_sll_482_M1_2_35 ( .A(u4_sll_482_ML_int_2__35_), .B(
        u4_sll_482_ML_int_2__31_), .S(u4_sll_482_n28), .Z(
        u4_sll_482_ML_int_3__35_) );
  MUX2_X2 u4_sll_482_M1_2_36 ( .A(u4_sll_482_ML_int_2__36_), .B(
        u4_sll_482_ML_int_2__32_), .S(u4_sll_482_n29), .Z(
        u4_sll_482_ML_int_3__36_) );
  MUX2_X2 u4_sll_482_M1_2_37 ( .A(u4_sll_482_ML_int_2__37_), .B(
        u4_sll_482_ML_int_2__33_), .S(u4_sll_482_n25), .Z(
        u4_sll_482_ML_int_3__37_) );
  MUX2_X2 u4_sll_482_M1_2_38 ( .A(u4_sll_482_ML_int_2__38_), .B(
        u4_sll_482_ML_int_2__34_), .S(u4_sll_482_n25), .Z(
        u4_sll_482_ML_int_3__38_) );
  MUX2_X2 u4_sll_482_M1_2_39 ( .A(u4_sll_482_ML_int_2__39_), .B(
        u4_sll_482_ML_int_2__35_), .S(u4_sll_482_n25), .Z(
        u4_sll_482_ML_int_3__39_) );
  MUX2_X2 u4_sll_482_M1_2_40 ( .A(u4_sll_482_ML_int_2__40_), .B(
        u4_sll_482_ML_int_2__36_), .S(u4_sll_482_n25), .Z(
        u4_sll_482_ML_int_3__40_) );
  MUX2_X2 u4_sll_482_M1_2_41 ( .A(u4_sll_482_ML_int_2__41_), .B(
        u4_sll_482_ML_int_2__37_), .S(u4_sll_482_n25), .Z(
        u4_sll_482_ML_int_3__41_) );
  MUX2_X2 u4_sll_482_M1_2_42 ( .A(u4_sll_482_ML_int_2__42_), .B(
        u4_sll_482_ML_int_2__38_), .S(u4_sll_482_n25), .Z(
        u4_sll_482_ML_int_3__42_) );
  MUX2_X2 u4_sll_482_M1_2_43 ( .A(u4_sll_482_ML_int_2__43_), .B(
        u4_sll_482_ML_int_2__39_), .S(u4_sll_482_n25), .Z(
        u4_sll_482_ML_int_3__43_) );
  MUX2_X2 u4_sll_482_M1_2_44 ( .A(u4_sll_482_ML_int_2__44_), .B(
        u4_sll_482_ML_int_2__40_), .S(u4_sll_482_n25), .Z(
        u4_sll_482_ML_int_3__44_) );
  MUX2_X2 u4_sll_482_M1_2_45 ( .A(u4_sll_482_ML_int_2__45_), .B(
        u4_sll_482_ML_int_2__41_), .S(u4_sll_482_n25), .Z(
        u4_sll_482_ML_int_3__45_) );
  MUX2_X2 u4_sll_482_M1_2_46 ( .A(u4_sll_482_ML_int_2__46_), .B(
        u4_sll_482_ML_int_2__42_), .S(u4_sll_482_n25), .Z(
        u4_sll_482_ML_int_3__46_) );
  MUX2_X2 u4_sll_482_M1_2_47 ( .A(u4_sll_482_ML_int_2__47_), .B(
        u4_sll_482_ML_int_2__43_), .S(u4_sll_482_n25), .Z(
        u4_sll_482_ML_int_3__47_) );
  MUX2_X2 u4_sll_482_M1_2_48 ( .A(u4_sll_482_ML_int_2__48_), .B(
        u4_sll_482_ML_int_2__44_), .S(u4_sll_482_n26), .Z(
        u4_sll_482_ML_int_3__48_) );
  MUX2_X2 u4_sll_482_M1_2_49 ( .A(u4_sll_482_ML_int_2__49_), .B(
        u4_sll_482_ML_int_2__45_), .S(u4_sll_482_n26), .Z(
        u4_sll_482_ML_int_3__49_) );
  MUX2_X2 u4_sll_482_M1_2_50 ( .A(u4_sll_482_ML_int_2__50_), .B(
        u4_sll_482_ML_int_2__46_), .S(u4_sll_482_n26), .Z(
        u4_sll_482_ML_int_3__50_) );
  MUX2_X2 u4_sll_482_M1_2_51 ( .A(u4_sll_482_ML_int_2__51_), .B(
        u4_sll_482_ML_int_2__47_), .S(u4_sll_482_n26), .Z(
        u4_sll_482_ML_int_3__51_) );
  MUX2_X2 u4_sll_482_M1_2_52 ( .A(u4_sll_482_ML_int_2__52_), .B(
        u4_sll_482_ML_int_2__48_), .S(u4_sll_482_n26), .Z(
        u4_sll_482_ML_int_3__52_) );
  MUX2_X2 u4_sll_482_M1_2_53 ( .A(u4_sll_482_ML_int_2__53_), .B(
        u4_sll_482_ML_int_2__49_), .S(u4_sll_482_n26), .Z(
        u4_sll_482_ML_int_3__53_) );
  MUX2_X2 u4_sll_482_M1_2_54 ( .A(u4_sll_482_ML_int_2__54_), .B(
        u4_sll_482_ML_int_2__50_), .S(u4_sll_482_n26), .Z(
        u4_sll_482_ML_int_3__54_) );
  MUX2_X2 u4_sll_482_M1_2_55 ( .A(u4_sll_482_ML_int_2__55_), .B(
        u4_sll_482_ML_int_2__51_), .S(u4_sll_482_n26), .Z(
        u4_sll_482_ML_int_3__55_) );
  MUX2_X2 u4_sll_482_M1_2_56 ( .A(u4_sll_482_ML_int_2__56_), .B(
        u4_sll_482_ML_int_2__52_), .S(u4_sll_482_n26), .Z(
        u4_sll_482_ML_int_3__56_) );
  MUX2_X2 u4_sll_482_M1_2_57 ( .A(u4_sll_482_ML_int_2__57_), .B(
        u4_sll_482_ML_int_2__53_), .S(u4_sll_482_n26), .Z(
        u4_sll_482_ML_int_3__57_) );
  MUX2_X2 u4_sll_482_M1_2_58 ( .A(u4_sll_482_ML_int_2__58_), .B(
        u4_sll_482_ML_int_2__54_), .S(u4_sll_482_n26), .Z(
        u4_sll_482_ML_int_3__58_) );
  MUX2_X2 u4_sll_482_M1_2_59 ( .A(u4_sll_482_ML_int_2__59_), .B(
        u4_sll_482_ML_int_2__55_), .S(u4_sll_482_n28), .Z(
        u4_sll_482_ML_int_3__59_) );
  MUX2_X2 u4_sll_482_M1_2_60 ( .A(u4_sll_482_ML_int_2__60_), .B(
        u4_sll_482_ML_int_2__56_), .S(u4_sll_482_n26), .Z(
        u4_sll_482_ML_int_3__60_) );
  MUX2_X2 u4_sll_482_M1_2_61 ( .A(u4_sll_482_ML_int_2__61_), .B(
        u4_sll_482_ML_int_2__57_), .S(u4_sll_482_n28), .Z(
        u4_sll_482_ML_int_3__61_) );
  MUX2_X2 u4_sll_482_M1_2_62 ( .A(u4_sll_482_ML_int_2__62_), .B(
        u4_sll_482_ML_int_2__58_), .S(u4_sll_482_n25), .Z(
        u4_sll_482_ML_int_3__62_) );
  MUX2_X2 u4_sll_482_M1_2_63 ( .A(u4_sll_482_ML_int_2__63_), .B(
        u4_sll_482_ML_int_2__59_), .S(u4_sll_482_n26), .Z(
        u4_sll_482_ML_int_3__63_) );
  MUX2_X2 u4_sll_482_M1_2_64 ( .A(u4_sll_482_ML_int_2__64_), .B(
        u4_sll_482_ML_int_2__60_), .S(u4_sll_482_n28), .Z(
        u4_sll_482_ML_int_3__64_) );
  MUX2_X2 u4_sll_482_M1_2_65 ( .A(u4_sll_482_ML_int_2__65_), .B(
        u4_sll_482_ML_int_2__61_), .S(u4_sll_482_n25), .Z(
        u4_sll_482_ML_int_3__65_) );
  MUX2_X2 u4_sll_482_M1_2_66 ( .A(u4_sll_482_ML_int_2__66_), .B(
        u4_sll_482_ML_int_2__62_), .S(u4_sll_482_n25), .Z(
        u4_sll_482_ML_int_3__66_) );
  MUX2_X2 u4_sll_482_M1_2_67 ( .A(u4_sll_482_ML_int_2__67_), .B(
        u4_sll_482_ML_int_2__63_), .S(u4_sll_482_n28), .Z(
        u4_sll_482_ML_int_3__67_) );
  MUX2_X2 u4_sll_482_M1_2_68 ( .A(u4_sll_482_ML_int_2__68_), .B(
        u4_sll_482_ML_int_2__64_), .S(u4_sll_482_n23), .Z(
        u4_sll_482_ML_int_3__68_) );
  MUX2_X2 u4_sll_482_M1_2_69 ( .A(u4_sll_482_ML_int_2__69_), .B(
        u4_sll_482_ML_int_2__65_), .S(u4_sll_482_n24), .Z(
        u4_sll_482_ML_int_3__69_) );
  MUX2_X2 u4_sll_482_M1_2_70 ( .A(u4_sll_482_ML_int_2__70_), .B(
        u4_sll_482_ML_int_2__66_), .S(u4_sll_482_n27), .Z(
        u4_sll_482_ML_int_3__70_) );
  MUX2_X2 u4_sll_482_M1_2_71 ( .A(u4_sll_482_ML_int_2__71_), .B(
        u4_sll_482_ML_int_2__67_), .S(u4_sll_482_n27), .Z(
        u4_sll_482_ML_int_3__71_) );
  MUX2_X2 u4_sll_482_M1_2_72 ( .A(u4_sll_482_ML_int_2__72_), .B(
        u4_sll_482_ML_int_2__68_), .S(u4_sll_482_n27), .Z(
        u4_sll_482_ML_int_3__72_) );
  MUX2_X2 u4_sll_482_M1_2_73 ( .A(u4_sll_482_ML_int_2__73_), .B(
        u4_sll_482_ML_int_2__69_), .S(u4_sll_482_n27), .Z(
        u4_sll_482_ML_int_3__73_) );
  MUX2_X2 u4_sll_482_M1_2_74 ( .A(u4_sll_482_ML_int_2__74_), .B(
        u4_sll_482_ML_int_2__70_), .S(u4_sll_482_n27), .Z(
        u4_sll_482_ML_int_3__74_) );
  MUX2_X2 u4_sll_482_M1_2_75 ( .A(u4_sll_482_ML_int_2__75_), .B(
        u4_sll_482_ML_int_2__71_), .S(u4_sll_482_n27), .Z(
        u4_sll_482_ML_int_3__75_) );
  MUX2_X2 u4_sll_482_M1_2_76 ( .A(u4_sll_482_ML_int_2__76_), .B(
        u4_sll_482_ML_int_2__72_), .S(u4_sll_482_n27), .Z(
        u4_sll_482_ML_int_3__76_) );
  MUX2_X2 u4_sll_482_M1_2_77 ( .A(u4_sll_482_ML_int_2__77_), .B(
        u4_sll_482_ML_int_2__73_), .S(u4_sll_482_n27), .Z(
        u4_sll_482_ML_int_3__77_) );
  MUX2_X2 u4_sll_482_M1_2_78 ( .A(u4_sll_482_ML_int_2__78_), .B(
        u4_sll_482_ML_int_2__74_), .S(u4_sll_482_n27), .Z(
        u4_sll_482_ML_int_3__78_) );
  MUX2_X2 u4_sll_482_M1_2_79 ( .A(u4_sll_482_ML_int_2__79_), .B(
        u4_sll_482_ML_int_2__75_), .S(u4_sll_482_n27), .Z(
        u4_sll_482_ML_int_3__79_) );
  MUX2_X2 u4_sll_482_M1_2_80 ( .A(u4_sll_482_ML_int_2__80_), .B(
        u4_sll_482_ML_int_2__76_), .S(u4_sll_482_n27), .Z(
        u4_sll_482_ML_int_3__80_) );
  MUX2_X2 u4_sll_482_M1_2_81 ( .A(u4_sll_482_ML_int_2__81_), .B(
        u4_sll_482_ML_int_2__77_), .S(u4_sll_482_n27), .Z(
        u4_sll_482_ML_int_3__81_) );
  MUX2_X2 u4_sll_482_M1_2_82 ( .A(u4_sll_482_ML_int_2__82_), .B(
        u4_sll_482_ML_int_2__78_), .S(u4_sll_482_n27), .Z(
        u4_sll_482_ML_int_3__82_) );
  MUX2_X2 u4_sll_482_M1_2_83 ( .A(u4_sll_482_ML_int_2__83_), .B(
        u4_sll_482_ML_int_2__79_), .S(u4_sll_482_n27), .Z(
        u4_sll_482_ML_int_3__83_) );
  MUX2_X2 u4_sll_482_M1_2_84 ( .A(u4_sll_482_ML_int_2__84_), .B(
        u4_sll_482_ML_int_2__80_), .S(u4_sll_482_n27), .Z(
        u4_sll_482_ML_int_3__84_) );
  MUX2_X2 u4_sll_482_M1_2_85 ( .A(u4_sll_482_ML_int_2__85_), .B(
        u4_sll_482_ML_int_2__81_), .S(u4_sll_482_n27), .Z(
        u4_sll_482_ML_int_3__85_) );
  MUX2_X2 u4_sll_482_M1_2_86 ( .A(u4_sll_482_ML_int_2__86_), .B(
        u4_sll_482_ML_int_2__82_), .S(u4_sll_482_n27), .Z(
        u4_sll_482_ML_int_3__86_) );
  MUX2_X2 u4_sll_482_M1_2_87 ( .A(u4_sll_482_ML_int_2__87_), .B(
        u4_sll_482_ML_int_2__83_), .S(u4_sll_482_n27), .Z(
        u4_sll_482_ML_int_3__87_) );
  MUX2_X2 u4_sll_482_M1_2_88 ( .A(u4_sll_482_ML_int_2__88_), .B(
        u4_sll_482_ML_int_2__84_), .S(u4_sll_482_n27), .Z(
        u4_sll_482_ML_int_3__88_) );
  MUX2_X2 u4_sll_482_M1_2_89 ( .A(u4_sll_482_ML_int_2__89_), .B(
        u4_sll_482_ML_int_2__85_), .S(u4_sll_482_n27), .Z(
        u4_sll_482_ML_int_3__89_) );
  MUX2_X2 u4_sll_482_M1_2_90 ( .A(u4_sll_482_ML_int_2__90_), .B(
        u4_sll_482_ML_int_2__86_), .S(u4_sll_482_n27), .Z(
        u4_sll_482_ML_int_3__90_) );
  MUX2_X2 u4_sll_482_M1_2_91 ( .A(u4_sll_482_ML_int_2__91_), .B(
        u4_sll_482_ML_int_2__87_), .S(u4_sll_482_n27), .Z(
        u4_sll_482_ML_int_3__91_) );
  MUX2_X2 u4_sll_482_M1_2_92 ( .A(u4_sll_482_ML_int_2__92_), .B(
        u4_sll_482_ML_int_2__88_), .S(u4_sll_482_n28), .Z(
        u4_sll_482_ML_int_3__92_) );
  MUX2_X2 u4_sll_482_M1_2_93 ( .A(u4_sll_482_ML_int_2__93_), .B(
        u4_sll_482_ML_int_2__89_), .S(u4_sll_482_n28), .Z(
        u4_sll_482_ML_int_3__93_) );
  MUX2_X2 u4_sll_482_M1_2_94 ( .A(u4_sll_482_ML_int_2__94_), .B(
        u4_sll_482_ML_int_2__90_), .S(u4_sll_482_n28), .Z(
        u4_sll_482_ML_int_3__94_) );
  MUX2_X2 u4_sll_482_M1_2_95 ( .A(u4_sll_482_ML_int_2__95_), .B(
        u4_sll_482_ML_int_2__91_), .S(u4_sll_482_n28), .Z(
        u4_sll_482_ML_int_3__95_) );
  MUX2_X2 u4_sll_482_M1_2_96 ( .A(u4_sll_482_ML_int_2__96_), .B(
        u4_sll_482_ML_int_2__92_), .S(u4_sll_482_n28), .Z(
        u4_sll_482_ML_int_3__96_) );
  MUX2_X2 u4_sll_482_M1_2_97 ( .A(u4_sll_482_ML_int_2__97_), .B(
        u4_sll_482_ML_int_2__93_), .S(u4_sll_482_n28), .Z(
        u4_sll_482_ML_int_3__97_) );
  MUX2_X2 u4_sll_482_M1_2_98 ( .A(u4_sll_482_ML_int_2__98_), .B(
        u4_sll_482_ML_int_2__94_), .S(u4_sll_482_n28), .Z(
        u4_sll_482_ML_int_3__98_) );
  MUX2_X2 u4_sll_482_M1_2_99 ( .A(u4_sll_482_ML_int_2__99_), .B(
        u4_sll_482_ML_int_2__95_), .S(u4_sll_482_n28), .Z(
        u4_sll_482_ML_int_3__99_) );
  MUX2_X2 u4_sll_482_M1_2_100 ( .A(u4_sll_482_ML_int_2__100_), .B(
        u4_sll_482_ML_int_2__96_), .S(u4_sll_482_n28), .Z(
        u4_sll_482_ML_int_3__100_) );
  MUX2_X2 u4_sll_482_M1_2_101 ( .A(u4_sll_482_ML_int_2__101_), .B(
        u4_sll_482_ML_int_2__97_), .S(u4_sll_482_n28), .Z(
        u4_sll_482_ML_int_3__101_) );
  MUX2_X2 u4_sll_482_M1_2_102 ( .A(u4_sll_482_ML_int_2__102_), .B(
        u4_sll_482_ML_int_2__98_), .S(u4_sll_482_n28), .Z(
        u4_sll_482_ML_int_3__102_) );
  MUX2_X2 u4_sll_482_M1_2_103 ( .A(u4_sll_482_ML_int_2__103_), .B(
        u4_sll_482_ML_int_2__99_), .S(u4_sll_482_n29), .Z(
        u4_sll_482_ML_int_3__103_) );
  MUX2_X2 u4_sll_482_M1_2_104 ( .A(u4_sll_482_ML_int_2__104_), .B(
        u4_sll_482_ML_int_2__100_), .S(u4_sll_482_n29), .Z(
        u4_sll_482_ML_int_3__104_) );
  MUX2_X2 u4_sll_482_M1_2_105 ( .A(u4_sll_482_ML_int_2__105_), .B(
        u4_sll_482_ML_int_2__101_), .S(u4_sll_482_n29), .Z(
        u4_sll_482_ML_int_3__105_) );
  MUX2_X2 u4_sll_482_M1_2_106 ( .A(u4_sll_482_ML_int_2__106_), .B(
        u4_sll_482_ML_int_2__102_), .S(u4_sll_482_n29), .Z(
        u4_sll_482_ML_int_3__106_) );
  MUX2_X2 u4_sll_482_M1_2_107 ( .A(u4_sll_482_ML_int_2__107_), .B(
        u4_sll_482_ML_int_2__103_), .S(u4_sll_482_n29), .Z(
        u4_sll_482_ML_int_3__107_) );
  MUX2_X2 u4_sll_482_M1_2_108 ( .A(u4_sll_482_ML_int_2__108_), .B(
        u4_sll_482_ML_int_2__104_), .S(u4_sll_482_n29), .Z(
        u4_sll_482_ML_int_3__108_) );
  MUX2_X2 u4_sll_482_M1_2_109 ( .A(u4_sll_482_ML_int_2__109_), .B(
        u4_sll_482_ML_int_2__105_), .S(u4_sll_482_n29), .Z(
        u4_sll_482_ML_int_3__109_) );
  MUX2_X2 u4_sll_482_M1_2_110 ( .A(u4_sll_482_ML_int_2__110_), .B(
        u4_sll_482_ML_int_2__106_), .S(u4_sll_482_n29), .Z(
        u4_sll_482_ML_int_3__110_) );
  MUX2_X2 u4_sll_482_M1_2_111 ( .A(u4_sll_482_ML_int_2__111_), .B(
        u4_sll_482_ML_int_2__107_), .S(u4_sll_482_n29), .Z(
        u4_sll_482_ML_int_3__111_) );
  MUX2_X2 u4_sll_482_M1_2_112 ( .A(u4_sll_482_ML_int_2__112_), .B(
        u4_sll_482_ML_int_2__108_), .S(u4_sll_482_n29), .Z(
        u4_sll_482_ML_int_3__112_) );
  MUX2_X2 u4_sll_482_M1_2_113 ( .A(u4_sll_482_ML_int_2__113_), .B(
        u4_sll_482_ML_int_2__109_), .S(u4_sll_482_n29), .Z(
        u4_sll_482_ML_int_3__113_) );
  MUX2_X2 u4_sll_482_M1_2_114 ( .A(u4_sll_482_ML_int_2__114_), .B(
        u4_sll_482_ML_int_2__110_), .S(u4_sll_482_n29), .Z(
        u4_sll_482_ML_int_3__114_) );
  MUX2_X2 u4_sll_482_M1_2_115 ( .A(u4_sll_482_n3), .B(
        u4_sll_482_ML_int_2__111_), .S(u4_sll_482_n29), .Z(
        u4_sll_482_ML_int_3__115_) );
  MUX2_X2 u4_sll_482_M1_2_116 ( .A(u4_sll_482_n4), .B(
        u4_sll_482_ML_int_2__112_), .S(u4_sll_482_n29), .Z(
        u4_sll_482_ML_int_3__116_) );
  MUX2_X2 u4_sll_482_M1_3_11 ( .A(u4_sll_482_ML_int_3__11_), .B(u4_sll_482_n40), .S(u4_sll_482_n32), .Z(u4_sll_482_ML_int_4__11_) );
  MUX2_X2 u4_sll_482_M1_3_12 ( .A(u4_sll_482_ML_int_3__12_), .B(
        u4_sll_482_ML_int_3__4_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__12_) );
  MUX2_X2 u4_sll_482_M1_3_13 ( .A(u4_sll_482_ML_int_3__13_), .B(
        u4_sll_482_ML_int_3__5_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__13_) );
  MUX2_X2 u4_sll_482_M1_3_14 ( .A(u4_sll_482_ML_int_3__14_), .B(
        u4_sll_482_ML_int_3__6_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__14_) );
  MUX2_X2 u4_sll_482_M1_3_15 ( .A(u4_sll_482_ML_int_3__15_), .B(
        u4_sll_482_ML_int_3__7_), .S(u4_sll_482_temp_int_SH_3_), .Z(
        u4_sll_482_ML_int_4__15_) );
  MUX2_X2 u4_sll_482_M1_3_16 ( .A(u4_sll_482_ML_int_3__16_), .B(
        u4_sll_482_ML_int_3__8_), .S(u4_sll_482_temp_int_SH_3_), .Z(
        u4_sll_482_ML_int_4__16_) );
  MUX2_X2 u4_sll_482_M1_3_17 ( .A(u4_sll_482_ML_int_3__17_), .B(
        u4_sll_482_ML_int_3__9_), .S(u4_sll_482_temp_int_SH_3_), .Z(
        u4_sll_482_ML_int_4__17_) );
  MUX2_X2 u4_sll_482_M1_3_18 ( .A(u4_sll_482_ML_int_3__18_), .B(
        u4_sll_482_ML_int_3__10_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__18_) );
  MUX2_X2 u4_sll_482_M1_3_19 ( .A(u4_sll_482_ML_int_3__19_), .B(
        u4_sll_482_ML_int_3__11_), .S(u4_sll_482_n30), .Z(
        u4_sll_482_ML_int_4__19_) );
  MUX2_X2 u4_sll_482_M1_3_20 ( .A(u4_sll_482_ML_int_3__20_), .B(
        u4_sll_482_ML_int_3__12_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__20_) );
  MUX2_X2 u4_sll_482_M1_3_21 ( .A(u4_sll_482_ML_int_3__21_), .B(
        u4_sll_482_ML_int_3__13_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__21_) );
  MUX2_X2 u4_sll_482_M1_3_27 ( .A(u4_sll_482_ML_int_3__27_), .B(
        u4_sll_482_ML_int_3__19_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__27_) );
  MUX2_X2 u4_sll_482_M1_3_28 ( .A(u4_sll_482_ML_int_3__28_), .B(
        u4_sll_482_ML_int_3__20_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__28_) );
  MUX2_X2 u4_sll_482_M1_3_29 ( .A(u4_sll_482_ML_int_3__29_), .B(
        u4_sll_482_ML_int_3__21_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__29_) );
  MUX2_X2 u4_sll_482_M1_3_30 ( .A(u4_sll_482_ML_int_3__30_), .B(
        u4_sll_482_ML_int_3__22_), .S(u4_sll_482_temp_int_SH_3_), .Z(
        u4_sll_482_ML_int_4__30_) );
  MUX2_X2 u4_sll_482_M1_3_31 ( .A(u4_sll_482_ML_int_3__31_), .B(
        u4_sll_482_ML_int_3__23_), .S(u4_sll_482_temp_int_SH_3_), .Z(
        u4_sll_482_ML_int_4__31_) );
  MUX2_X2 u4_sll_482_M1_3_32 ( .A(u4_sll_482_ML_int_3__32_), .B(
        u4_sll_482_ML_int_3__24_), .S(u4_sll_482_temp_int_SH_3_), .Z(
        u4_sll_482_ML_int_4__32_) );
  MUX2_X2 u4_sll_482_M1_3_33 ( .A(u4_sll_482_ML_int_3__33_), .B(
        u4_sll_482_ML_int_3__25_), .S(u4_sll_482_temp_int_SH_3_), .Z(
        u4_sll_482_ML_int_4__33_) );
  MUX2_X2 u4_sll_482_M1_3_34 ( .A(u4_sll_482_ML_int_3__34_), .B(
        u4_sll_482_ML_int_3__26_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__34_) );
  MUX2_X2 u4_sll_482_M1_3_35 ( .A(u4_sll_482_ML_int_3__35_), .B(
        u4_sll_482_ML_int_3__27_), .S(u4_sll_482_n30), .Z(
        u4_sll_482_ML_int_4__35_) );
  MUX2_X2 u4_sll_482_M1_3_36 ( .A(u4_sll_482_ML_int_3__36_), .B(
        u4_sll_482_ML_int_3__28_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__36_) );
  MUX2_X2 u4_sll_482_M1_3_37 ( .A(u4_sll_482_ML_int_3__37_), .B(
        u4_sll_482_ML_int_3__29_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__37_) );
  MUX2_X2 u4_sll_482_M1_3_43 ( .A(u4_sll_482_ML_int_3__43_), .B(
        u4_sll_482_ML_int_3__35_), .S(u4_sll_482_n31), .Z(
        u4_sll_482_ML_int_4__43_) );
  MUX2_X2 u4_sll_482_M1_3_44 ( .A(u4_sll_482_ML_int_3__44_), .B(
        u4_sll_482_ML_int_3__36_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__44_) );
  MUX2_X2 u4_sll_482_M1_3_45 ( .A(u4_sll_482_ML_int_3__45_), .B(
        u4_sll_482_ML_int_3__37_), .S(u4_sll_482_n31), .Z(
        u4_sll_482_ML_int_4__45_) );
  MUX2_X2 u4_sll_482_M1_3_46 ( .A(u4_sll_482_ML_int_3__46_), .B(
        u4_sll_482_ML_int_3__38_), .S(u4_sll_482_temp_int_SH_3_), .Z(
        u4_sll_482_ML_int_4__46_) );
  MUX2_X2 u4_sll_482_M1_3_47 ( .A(u4_sll_482_ML_int_3__47_), .B(
        u4_sll_482_ML_int_3__39_), .S(u4_sll_482_n30), .Z(
        u4_sll_482_ML_int_4__47_) );
  MUX2_X2 u4_sll_482_M1_3_48 ( .A(u4_sll_482_ML_int_3__48_), .B(
        u4_sll_482_ML_int_3__40_), .S(u4_sll_482_temp_int_SH_3_), .Z(
        u4_sll_482_ML_int_4__48_) );
  MUX2_X2 u4_sll_482_M1_3_49 ( .A(u4_sll_482_ML_int_3__49_), .B(
        u4_sll_482_ML_int_3__41_), .S(u4_sll_482_n30), .Z(
        u4_sll_482_ML_int_4__49_) );
  MUX2_X2 u4_sll_482_M1_3_50 ( .A(u4_sll_482_ML_int_3__50_), .B(
        u4_sll_482_ML_int_3__42_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__50_) );
  MUX2_X2 u4_sll_482_M1_3_51 ( .A(u4_sll_482_ML_int_3__51_), .B(
        u4_sll_482_ML_int_3__43_), .S(u4_sll_482_n31), .Z(
        u4_sll_482_ML_int_4__51_) );
  MUX2_X2 u4_sll_482_M1_3_52 ( .A(u4_sll_482_ML_int_3__52_), .B(
        u4_sll_482_ML_int_3__44_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__52_) );
  MUX2_X2 u4_sll_482_M1_3_53 ( .A(u4_sll_482_ML_int_3__53_), .B(
        u4_sll_482_ML_int_3__45_), .S(u4_sll_482_n31), .Z(
        u4_sll_482_ML_int_4__53_) );
  MUX2_X2 u4_sll_482_M1_3_59 ( .A(u4_sll_482_ML_int_3__59_), .B(
        u4_sll_482_ML_int_3__51_), .S(u4_sll_482_n31), .Z(
        u4_sll_482_ML_int_4__59_) );
  MUX2_X2 u4_sll_482_M1_3_60 ( .A(u4_sll_482_ML_int_3__60_), .B(
        u4_sll_482_ML_int_3__52_), .S(u4_sll_482_n31), .Z(
        u4_sll_482_ML_int_4__60_) );
  MUX2_X2 u4_sll_482_M1_3_61 ( .A(u4_sll_482_ML_int_3__61_), .B(
        u4_sll_482_ML_int_3__53_), .S(u4_sll_482_n31), .Z(
        u4_sll_482_ML_int_4__61_) );
  MUX2_X2 u4_sll_482_M1_3_62 ( .A(u4_sll_482_ML_int_3__62_), .B(
        u4_sll_482_ML_int_3__54_), .S(u4_sll_482_n31), .Z(
        u4_sll_482_ML_int_4__62_) );
  MUX2_X2 u4_sll_482_M1_3_63 ( .A(u4_sll_482_ML_int_3__63_), .B(
        u4_sll_482_ML_int_3__55_), .S(u4_sll_482_n31), .Z(
        u4_sll_482_ML_int_4__63_) );
  MUX2_X2 u4_sll_482_M1_3_64 ( .A(u4_sll_482_ML_int_3__64_), .B(
        u4_sll_482_ML_int_3__56_), .S(u4_sll_482_n31), .Z(
        u4_sll_482_ML_int_4__64_) );
  MUX2_X2 u4_sll_482_M1_3_65 ( .A(u4_sll_482_ML_int_3__65_), .B(
        u4_sll_482_ML_int_3__57_), .S(u4_sll_482_n31), .Z(
        u4_sll_482_ML_int_4__65_) );
  MUX2_X2 u4_sll_482_M1_3_66 ( .A(u4_sll_482_ML_int_3__66_), .B(
        u4_sll_482_ML_int_3__58_), .S(u4_sll_482_n31), .Z(
        u4_sll_482_ML_int_4__66_) );
  MUX2_X2 u4_sll_482_M1_3_67 ( .A(u4_sll_482_ML_int_3__67_), .B(
        u4_sll_482_ML_int_3__59_), .S(u4_sll_482_n31), .Z(
        u4_sll_482_ML_int_4__67_) );
  MUX2_X2 u4_sll_482_M1_3_68 ( .A(u4_sll_482_ML_int_3__68_), .B(
        u4_sll_482_ML_int_3__60_), .S(u4_sll_482_n31), .Z(
        u4_sll_482_ML_int_4__68_) );
  MUX2_X2 u4_sll_482_M1_3_69 ( .A(u4_sll_482_ML_int_3__69_), .B(
        u4_sll_482_ML_int_3__61_), .S(u4_sll_482_n31), .Z(
        u4_sll_482_ML_int_4__69_) );
  MUX2_X2 u4_sll_482_M1_3_75 ( .A(u4_sll_482_ML_int_3__75_), .B(
        u4_sll_482_ML_int_3__67_), .S(u4_sll_482_n30), .Z(
        u4_sll_482_ML_int_4__75_) );
  MUX2_X2 u4_sll_482_M1_3_76 ( .A(u4_sll_482_ML_int_3__76_), .B(
        u4_sll_482_ML_int_3__68_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__76_) );
  MUX2_X2 u4_sll_482_M1_3_77 ( .A(u4_sll_482_ML_int_3__77_), .B(
        u4_sll_482_ML_int_3__69_), .S(u4_sll_482_n30), .Z(
        u4_sll_482_ML_int_4__77_) );
  MUX2_X2 u4_sll_482_M1_3_78 ( .A(u4_sll_482_ML_int_3__78_), .B(
        u4_sll_482_ML_int_3__70_), .S(u4_sll_482_temp_int_SH_3_), .Z(
        u4_sll_482_ML_int_4__78_) );
  MUX2_X2 u4_sll_482_M1_3_79 ( .A(u4_sll_482_ML_int_3__79_), .B(
        u4_sll_482_ML_int_3__71_), .S(u4_sll_482_n31), .Z(
        u4_sll_482_ML_int_4__79_) );
  MUX2_X2 u4_sll_482_M1_3_80 ( .A(u4_sll_482_ML_int_3__80_), .B(
        u4_sll_482_ML_int_3__72_), .S(u4_sll_482_temp_int_SH_3_), .Z(
        u4_sll_482_ML_int_4__80_) );
  MUX2_X2 u4_sll_482_M1_3_81 ( .A(u4_sll_482_ML_int_3__81_), .B(
        u4_sll_482_ML_int_3__73_), .S(u4_sll_482_n30), .Z(
        u4_sll_482_ML_int_4__81_) );
  MUX2_X2 u4_sll_482_M1_3_82 ( .A(u4_sll_482_ML_int_3__82_), .B(
        u4_sll_482_ML_int_3__74_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__82_) );
  MUX2_X2 u4_sll_482_M1_3_83 ( .A(u4_sll_482_ML_int_3__83_), .B(
        u4_sll_482_ML_int_3__75_), .S(u4_sll_482_temp_int_SH_3_), .Z(
        u4_sll_482_ML_int_4__83_) );
  MUX2_X2 u4_sll_482_M1_3_84 ( .A(u4_sll_482_ML_int_3__84_), .B(
        u4_sll_482_ML_int_3__76_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__84_) );
  MUX2_X2 u4_sll_482_M1_3_85 ( .A(u4_sll_482_ML_int_3__85_), .B(
        u4_sll_482_ML_int_3__77_), .S(u4_sll_482_n30), .Z(
        u4_sll_482_ML_int_4__85_) );
  MUX2_X2 u4_sll_482_M1_3_91 ( .A(u4_sll_482_ML_int_3__91_), .B(
        u4_sll_482_ML_int_3__83_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__91_) );
  MUX2_X2 u4_sll_482_M1_3_92 ( .A(u4_sll_482_ML_int_3__92_), .B(
        u4_sll_482_ML_int_3__84_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__92_) );
  MUX2_X2 u4_sll_482_M1_3_93 ( .A(u4_sll_482_ML_int_3__93_), .B(
        u4_sll_482_ML_int_3__85_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__93_) );
  MUX2_X2 u4_sll_482_M1_3_94 ( .A(u4_sll_482_ML_int_3__94_), .B(
        u4_sll_482_ML_int_3__86_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__94_) );
  MUX2_X2 u4_sll_482_M1_3_95 ( .A(u4_sll_482_ML_int_3__95_), .B(
        u4_sll_482_ML_int_3__87_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__95_) );
  MUX2_X2 u4_sll_482_M1_3_96 ( .A(u4_sll_482_ML_int_3__96_), .B(
        u4_sll_482_ML_int_3__88_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__96_) );
  MUX2_X2 u4_sll_482_M1_3_97 ( .A(u4_sll_482_ML_int_3__97_), .B(
        u4_sll_482_ML_int_3__89_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__97_) );
  MUX2_X2 u4_sll_482_M1_3_98 ( .A(u4_sll_482_ML_int_3__98_), .B(
        u4_sll_482_ML_int_3__90_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__98_) );
  MUX2_X2 u4_sll_482_M1_3_99 ( .A(u4_sll_482_ML_int_3__99_), .B(
        u4_sll_482_ML_int_3__91_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__99_) );
  MUX2_X2 u4_sll_482_M1_3_100 ( .A(u4_sll_482_ML_int_3__100_), .B(
        u4_sll_482_ML_int_3__92_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__100_) );
  MUX2_X2 u4_sll_482_M1_3_101 ( .A(u4_sll_482_ML_int_3__101_), .B(
        u4_sll_482_ML_int_3__93_), .S(u4_sll_482_n32), .Z(
        u4_sll_482_ML_int_4__101_) );
  MUX2_X2 u4_sll_482_M1_3_107 ( .A(u4_sll_482_ML_int_3__107_), .B(
        u4_sll_482_ML_int_3__99_), .S(u4_sll_482_n30), .Z(
        u4_sll_482_ML_int_4__107_) );
  MUX2_X2 u4_sll_482_M1_3_108 ( .A(u4_sll_482_ML_int_3__108_), .B(
        u4_sll_482_ML_int_3__100_), .S(u4_sll_482_n30), .Z(
        u4_sll_482_ML_int_4__108_) );
  MUX2_X2 u4_sll_482_M1_3_109 ( .A(u4_sll_482_ML_int_3__109_), .B(
        u4_sll_482_ML_int_3__101_), .S(u4_sll_482_n30), .Z(
        u4_sll_482_ML_int_4__109_) );
  MUX2_X2 u4_sll_482_M1_3_110 ( .A(u4_sll_482_ML_int_3__110_), .B(
        u4_sll_482_ML_int_3__102_), .S(u4_sll_482_n30), .Z(
        u4_sll_482_ML_int_4__110_) );
  MUX2_X2 u4_sll_482_M1_3_111 ( .A(u4_sll_482_ML_int_3__111_), .B(
        u4_sll_482_ML_int_3__103_), .S(u4_sll_482_n30), .Z(
        u4_sll_482_ML_int_4__111_) );
  MUX2_X2 u4_sll_482_M1_3_112 ( .A(u4_sll_482_ML_int_3__112_), .B(
        u4_sll_482_ML_int_3__104_), .S(u4_sll_482_n30), .Z(
        u4_sll_482_ML_int_4__112_) );
  MUX2_X2 u4_sll_482_M1_3_113 ( .A(u4_sll_482_ML_int_3__113_), .B(
        u4_sll_482_ML_int_3__105_), .S(u4_sll_482_n30), .Z(
        u4_sll_482_ML_int_4__113_) );
  MUX2_X2 u4_sll_482_M1_3_114 ( .A(u4_sll_482_ML_int_3__114_), .B(
        u4_sll_482_ML_int_3__106_), .S(u4_sll_482_n30), .Z(
        u4_sll_482_ML_int_4__114_) );
  MUX2_X2 u4_sll_482_M1_3_115 ( .A(u4_sll_482_ML_int_3__115_), .B(
        u4_sll_482_ML_int_3__107_), .S(u4_sll_482_n30), .Z(
        u4_sll_482_ML_int_4__115_) );
  MUX2_X2 u4_sll_482_M1_3_116 ( .A(u4_sll_482_ML_int_3__116_), .B(
        u4_sll_482_ML_int_3__108_), .S(u4_sll_482_n30), .Z(
        u4_sll_482_ML_int_4__116_) );
  MUX2_X2 u4_sll_482_M1_3_117 ( .A(u4_sll_482_n5), .B(
        u4_sll_482_ML_int_3__109_), .S(u4_sll_482_n30), .Z(
        u4_sll_482_ML_int_4__117_) );
  MUX2_X2 u4_sll_482_M1_4_16 ( .A(u4_sll_482_ML_int_4__16_), .B(
        u4_sll_482_ML_int_4__0_), .S(u4_sll_482_n35), .Z(
        u4_sll_482_ML_int_5__16_) );
  MUX2_X2 u4_sll_482_M1_4_17 ( .A(u4_sll_482_ML_int_4__17_), .B(
        u4_sll_482_ML_int_4__1_), .S(u4_sll_482_n35), .Z(
        u4_sll_482_ML_int_5__17_) );
  MUX2_X2 u4_sll_482_M1_4_18 ( .A(u4_sll_482_ML_int_4__18_), .B(
        u4_sll_482_ML_int_4__2_), .S(u4_sll_482_n36), .Z(
        u4_sll_482_ML_int_5__18_) );
  MUX2_X2 u4_sll_482_M1_4_19 ( .A(u4_sll_482_ML_int_4__19_), .B(
        u4_sll_482_ML_int_4__3_), .S(u4_sll_482_n35), .Z(
        u4_sll_482_ML_int_5__19_) );
  MUX2_X2 u4_sll_482_M1_4_20 ( .A(u4_sll_482_ML_int_4__20_), .B(
        u4_sll_482_ML_int_4__4_), .S(u4_sll_482_temp_int_SH_4_), .Z(
        u4_sll_482_ML_int_5__20_) );
  MUX2_X2 u4_sll_482_M1_4_21 ( .A(u4_sll_482_ML_int_4__21_), .B(
        u4_sll_482_ML_int_4__5_), .S(u4_sll_482_temp_int_SH_4_), .Z(
        u4_sll_482_ML_int_5__21_) );
  MUX2_X2 u4_sll_482_M1_4_43 ( .A(u4_sll_482_ML_int_4__43_), .B(
        u4_sll_482_ML_int_4__27_), .S(u4_sll_482_temp_int_SH_4_), .Z(
        u4_sll_482_ML_int_5__43_) );
  MUX2_X2 u4_sll_482_M1_4_44 ( .A(u4_sll_482_ML_int_4__44_), .B(
        u4_sll_482_ML_int_4__28_), .S(u4_sll_482_temp_int_SH_4_), .Z(
        u4_sll_482_ML_int_5__44_) );
  MUX2_X2 u4_sll_482_M1_4_45 ( .A(u4_sll_482_ML_int_4__45_), .B(
        u4_sll_482_ML_int_4__29_), .S(u4_sll_482_temp_int_SH_4_), .Z(
        u4_sll_482_ML_int_5__45_) );
  MUX2_X2 u4_sll_482_M1_4_46 ( .A(u4_sll_482_ML_int_4__46_), .B(
        u4_sll_482_ML_int_4__30_), .S(u4_sll_482_temp_int_SH_4_), .Z(
        u4_sll_482_ML_int_5__46_) );
  MUX2_X2 u4_sll_482_M1_4_47 ( .A(u4_sll_482_ML_int_4__47_), .B(
        u4_sll_482_ML_int_4__31_), .S(u4_sll_482_temp_int_SH_4_), .Z(
        u4_sll_482_ML_int_5__47_) );
  MUX2_X2 u4_sll_482_M1_4_48 ( .A(u4_sll_482_ML_int_4__48_), .B(
        u4_sll_482_ML_int_4__32_), .S(u4_sll_482_n35), .Z(
        u4_sll_482_ML_int_5__48_) );
  MUX2_X2 u4_sll_482_M1_4_49 ( .A(u4_sll_482_ML_int_4__49_), .B(
        u4_sll_482_ML_int_4__33_), .S(u4_sll_482_n35), .Z(
        u4_sll_482_ML_int_5__49_) );
  MUX2_X2 u4_sll_482_M1_4_50 ( .A(u4_sll_482_ML_int_4__50_), .B(
        u4_sll_482_ML_int_4__34_), .S(u4_sll_482_n35), .Z(
        u4_sll_482_ML_int_5__50_) );
  MUX2_X2 u4_sll_482_M1_4_51 ( .A(u4_sll_482_ML_int_4__51_), .B(
        u4_sll_482_ML_int_4__35_), .S(u4_sll_482_n35), .Z(
        u4_sll_482_ML_int_5__51_) );
  MUX2_X2 u4_sll_482_M1_4_52 ( .A(u4_sll_482_ML_int_4__52_), .B(
        u4_sll_482_ML_int_4__36_), .S(u4_sll_482_n35), .Z(
        u4_sll_482_ML_int_5__52_) );
  MUX2_X2 u4_sll_482_M1_4_53 ( .A(u4_sll_482_ML_int_4__53_), .B(
        u4_sll_482_ML_int_4__37_), .S(u4_sll_482_n35), .Z(
        u4_sll_482_ML_int_5__53_) );
  MUX2_X2 u4_sll_482_M1_4_75 ( .A(u4_sll_482_ML_int_4__75_), .B(
        u4_sll_482_ML_int_4__59_), .S(u4_sll_482_n35), .Z(
        u4_sll_482_ML_int_5__75_) );
  MUX2_X2 u4_sll_482_M1_4_76 ( .A(u4_sll_482_ML_int_4__76_), .B(
        u4_sll_482_ML_int_4__60_), .S(u4_sll_482_n35), .Z(
        u4_sll_482_ML_int_5__76_) );
  MUX2_X2 u4_sll_482_M1_4_77 ( .A(u4_sll_482_ML_int_4__77_), .B(
        u4_sll_482_ML_int_4__61_), .S(u4_sll_482_n35), .Z(
        u4_sll_482_ML_int_5__77_) );
  MUX2_X2 u4_sll_482_M1_4_78 ( .A(u4_sll_482_ML_int_4__78_), .B(
        u4_sll_482_ML_int_4__62_), .S(u4_sll_482_n35), .Z(
        u4_sll_482_ML_int_5__78_) );
  MUX2_X2 u4_sll_482_M1_4_79 ( .A(u4_sll_482_ML_int_4__79_), .B(
        u4_sll_482_ML_int_4__63_), .S(u4_sll_482_n35), .Z(
        u4_sll_482_ML_int_5__79_) );
  MUX2_X2 u4_sll_482_M1_4_80 ( .A(u4_sll_482_ML_int_4__80_), .B(
        u4_sll_482_ML_int_4__64_), .S(u4_sll_482_n36), .Z(
        u4_sll_482_ML_int_5__80_) );
  MUX2_X2 u4_sll_482_M1_4_81 ( .A(u4_sll_482_ML_int_4__81_), .B(
        u4_sll_482_ML_int_4__65_), .S(u4_sll_482_n36), .Z(
        u4_sll_482_ML_int_5__81_) );
  MUX2_X2 u4_sll_482_M1_4_82 ( .A(u4_sll_482_ML_int_4__82_), .B(
        u4_sll_482_ML_int_4__66_), .S(u4_sll_482_n36), .Z(
        u4_sll_482_ML_int_5__82_) );
  MUX2_X2 u4_sll_482_M1_4_83 ( .A(u4_sll_482_ML_int_4__83_), .B(
        u4_sll_482_ML_int_4__67_), .S(u4_sll_482_n36), .Z(
        u4_sll_482_ML_int_5__83_) );
  MUX2_X2 u4_sll_482_M1_4_84 ( .A(u4_sll_482_ML_int_4__84_), .B(
        u4_sll_482_ML_int_4__68_), .S(u4_sll_482_n36), .Z(
        u4_sll_482_ML_int_5__84_) );
  MUX2_X2 u4_sll_482_M1_4_85 ( .A(u4_sll_482_ML_int_4__85_), .B(
        u4_sll_482_ML_int_4__69_), .S(u4_sll_482_n36), .Z(
        u4_sll_482_ML_int_5__85_) );
  MUX2_X2 u4_sll_482_M1_4_107 ( .A(u4_sll_482_ML_int_4__107_), .B(
        u4_sll_482_ML_int_4__91_), .S(u4_sll_482_n36), .Z(
        u4_sll_482_ML_int_5__107_) );
  MUX2_X2 u4_sll_482_M1_4_108 ( .A(u4_sll_482_ML_int_4__108_), .B(
        u4_sll_482_ML_int_4__92_), .S(u4_sll_482_n36), .Z(
        u4_sll_482_ML_int_5__108_) );
  MUX2_X2 u4_sll_482_M1_4_109 ( .A(u4_sll_482_ML_int_4__109_), .B(
        u4_sll_482_ML_int_4__93_), .S(u4_sll_482_n36), .Z(
        u4_sll_482_ML_int_5__109_) );
  MUX2_X2 u4_sll_482_M1_4_110 ( .A(u4_sll_482_ML_int_4__110_), .B(
        u4_sll_482_ML_int_4__94_), .S(u4_sll_482_n36), .Z(
        u4_sll_482_ML_int_5__110_) );
  MUX2_X2 u4_sll_482_M1_4_111 ( .A(u4_sll_482_ML_int_4__111_), .B(
        u4_sll_482_ML_int_4__95_), .S(u4_sll_482_n36), .Z(
        u4_sll_482_ML_int_5__111_) );
  MUX2_X2 u4_sll_482_M1_4_112 ( .A(u4_sll_482_ML_int_4__112_), .B(
        u4_sll_482_ML_int_4__96_), .S(u4_sll_482_n36), .Z(
        u4_sll_482_ML_int_5__112_) );
  MUX2_X2 u4_sll_482_M1_4_113 ( .A(u4_sll_482_ML_int_4__113_), .B(
        u4_sll_482_ML_int_4__97_), .S(u4_sll_482_n35), .Z(
        u4_sll_482_ML_int_5__113_) );
  MUX2_X2 u4_sll_482_M1_4_114 ( .A(u4_sll_482_ML_int_4__114_), .B(
        u4_sll_482_ML_int_4__98_), .S(u4_sll_482_n35), .Z(
        u4_sll_482_ML_int_5__114_) );
  MUX2_X2 u4_sll_482_M1_4_115 ( .A(u4_sll_482_ML_int_4__115_), .B(
        u4_sll_482_ML_int_4__99_), .S(u4_sll_482_n36), .Z(
        u4_sll_482_ML_int_5__115_) );
  MUX2_X2 u4_sll_482_M1_4_116 ( .A(u4_sll_482_ML_int_4__116_), .B(
        u4_sll_482_ML_int_4__100_), .S(u4_sll_482_n35), .Z(
        u4_sll_482_ML_int_5__116_) );
  MUX2_X2 u4_sll_482_M1_4_117 ( .A(u4_sll_482_ML_int_4__117_), .B(
        u4_sll_482_ML_int_4__101_), .S(u4_sll_482_n36), .Z(
        u4_sll_482_ML_int_5__117_) );
  MUX2_X2 u4_sll_482_M1_5_43 ( .A(u4_sll_482_ML_int_5__43_), .B(
        u4_sll_482_ML_int_5__11_), .S(u4_sll_482_n41), .Z(
        u4_sll_482_ML_int_6__43_) );
  MUX2_X2 u4_sll_482_M1_5_44 ( .A(u4_sll_482_ML_int_5__44_), .B(
        u4_sll_482_ML_int_5__12_), .S(u4_sll_482_n41), .Z(
        u4_sll_482_ML_int_6__44_) );
  MUX2_X2 u4_sll_482_M1_5_45 ( .A(u4_sll_482_ML_int_5__45_), .B(
        u4_sll_482_ML_int_5__13_), .S(u4_sll_482_n41), .Z(
        u4_sll_482_ML_int_6__45_) );
  MUX2_X2 u4_sll_482_M1_5_46 ( .A(u4_sll_482_ML_int_5__46_), .B(
        u4_sll_482_ML_int_5__14_), .S(u4_sll_482_n41), .Z(
        u4_sll_482_ML_int_6__46_) );
  MUX2_X2 u4_sll_482_M1_5_47 ( .A(u4_sll_482_ML_int_5__47_), .B(
        u4_sll_482_ML_int_5__15_), .S(u4_sll_482_n41), .Z(
        u4_sll_482_ML_int_6__47_) );
  MUX2_X2 u4_sll_482_M1_5_48 ( .A(u4_sll_482_ML_int_5__48_), .B(
        u4_sll_482_ML_int_5__16_), .S(u4_sll_482_n41), .Z(
        u4_sll_482_ML_int_6__48_) );
  MUX2_X2 u4_sll_482_M1_5_49 ( .A(u4_sll_482_ML_int_5__49_), .B(
        u4_sll_482_ML_int_5__17_), .S(u4_sll_482_n41), .Z(
        u4_sll_482_ML_int_6__49_) );
  MUX2_X2 u4_sll_482_M1_5_50 ( .A(u4_sll_482_ML_int_5__50_), .B(
        u4_sll_482_ML_int_5__18_), .S(u4_sll_482_n41), .Z(
        u4_sll_482_ML_int_6__50_) );
  MUX2_X2 u4_sll_482_M1_5_51 ( .A(u4_sll_482_ML_int_5__51_), .B(
        u4_sll_482_ML_int_5__19_), .S(u4_sll_482_n41), .Z(
        u4_sll_482_ML_int_6__51_) );
  MUX2_X2 u4_sll_482_M1_5_52 ( .A(u4_sll_482_ML_int_5__52_), .B(
        u4_sll_482_ML_int_5__20_), .S(u4_sll_482_n41), .Z(
        u4_sll_482_ML_int_6__52_) );
  MUX2_X2 u4_sll_482_M1_5_53 ( .A(u4_sll_482_ML_int_5__53_), .B(
        u4_sll_482_ML_int_5__21_), .S(u4_sll_482_n41), .Z(
        u4_sll_482_ML_int_6__53_) );
  MUX2_X2 u4_sll_482_M1_5_107 ( .A(u4_sll_482_ML_int_5__107_), .B(
        u4_sll_482_ML_int_5__75_), .S(u4_sll_482_n41), .Z(
        u4_sll_482_ML_int_6__107_) );
  MUX2_X2 u4_sll_482_M1_5_108 ( .A(u4_sll_482_ML_int_5__108_), .B(
        u4_sll_482_ML_int_5__76_), .S(u4_sll_482_n41), .Z(
        u4_sll_482_ML_int_6__108_) );
  MUX2_X2 u4_sll_482_M1_5_109 ( .A(u4_sll_482_ML_int_5__109_), .B(
        u4_sll_482_ML_int_5__77_), .S(u4_sll_482_n41), .Z(
        u4_sll_482_ML_int_6__109_) );
  MUX2_X2 u4_sll_482_M1_5_110 ( .A(u4_sll_482_ML_int_5__110_), .B(
        u4_sll_482_ML_int_5__78_), .S(u4_sll_482_n41), .Z(
        u4_sll_482_ML_int_6__110_) );
  MUX2_X2 u4_sll_482_M1_5_111 ( .A(u4_sll_482_ML_int_5__111_), .B(
        u4_sll_482_ML_int_5__79_), .S(u4_sll_482_n41), .Z(
        u4_sll_482_ML_int_6__111_) );
  MUX2_X2 u4_sll_482_M1_5_112 ( .A(u4_sll_482_ML_int_5__112_), .B(
        u4_sll_482_ML_int_5__80_), .S(u4_sll_482_n41), .Z(
        u4_sll_482_ML_int_6__112_) );
  MUX2_X2 u4_sll_482_M1_5_113 ( .A(u4_sll_482_ML_int_5__113_), .B(
        u4_sll_482_ML_int_5__81_), .S(u4_sll_482_n41), .Z(
        u4_sll_482_ML_int_6__113_) );
  MUX2_X2 u4_sll_482_M1_5_114 ( .A(u4_sll_482_ML_int_5__114_), .B(
        u4_sll_482_ML_int_5__82_), .S(u4_sll_482_n41), .Z(
        u4_sll_482_ML_int_6__114_) );
  MUX2_X2 u4_sll_482_M1_5_115 ( .A(u4_sll_482_ML_int_5__115_), .B(
        u4_sll_482_ML_int_5__83_), .S(u4_sll_482_n41), .Z(
        u4_sll_482_ML_int_6__115_) );
  MUX2_X2 u4_sll_482_M1_5_116 ( .A(u4_sll_482_ML_int_5__116_), .B(
        u4_sll_482_ML_int_5__84_), .S(u4_sll_482_n41), .Z(
        u4_sll_482_ML_int_6__116_) );
  MUX2_X2 u4_sll_482_M1_5_117 ( .A(u4_sll_482_ML_int_5__117_), .B(
        u4_sll_482_ML_int_5__85_), .S(u4_sll_482_n41), .Z(
        u4_sll_482_ML_int_6__117_) );
  MUX2_X2 u4_sll_482_M1_6_107 ( .A(u4_sll_482_ML_int_6__107_), .B(
        u4_sll_482_ML_int_6__43_), .S(u4_sll_482_n42), .Z(
        u4_sll_482_ML_int_7__107_) );
  MUX2_X2 u4_sll_482_M1_6_108 ( .A(u4_sll_482_ML_int_6__108_), .B(
        u4_sll_482_ML_int_6__44_), .S(u4_sll_482_n42), .Z(
        u4_sll_482_ML_int_7__108_) );
  MUX2_X2 u4_sll_482_M1_6_109 ( .A(u4_sll_482_ML_int_6__109_), .B(
        u4_sll_482_ML_int_6__45_), .S(u4_sll_482_n42), .Z(
        u4_sll_482_ML_int_7__109_) );
  MUX2_X2 u4_sll_482_M1_6_110 ( .A(u4_sll_482_ML_int_6__110_), .B(
        u4_sll_482_ML_int_6__46_), .S(u4_sll_482_n42), .Z(
        u4_sll_482_ML_int_7__110_) );
  MUX2_X2 u4_sll_482_M1_6_111 ( .A(u4_sll_482_ML_int_6__111_), .B(
        u4_sll_482_ML_int_6__47_), .S(u4_sll_482_n42), .Z(
        u4_sll_482_ML_int_7__111_) );
  MUX2_X2 u4_sll_482_M1_6_112 ( .A(u4_sll_482_ML_int_6__112_), .B(
        u4_sll_482_ML_int_6__48_), .S(u4_sll_482_n42), .Z(
        u4_sll_482_ML_int_7__112_) );
  MUX2_X2 u4_sll_482_M1_6_113 ( .A(u4_sll_482_ML_int_6__113_), .B(
        u4_sll_482_ML_int_6__49_), .S(u4_sll_482_n42), .Z(
        u4_sll_482_ML_int_7__113_) );
  MUX2_X2 u4_sll_482_M1_6_114 ( .A(u4_sll_482_ML_int_6__114_), .B(
        u4_sll_482_ML_int_6__50_), .S(u4_sll_482_n42), .Z(
        u4_sll_482_ML_int_7__114_) );
  MUX2_X2 u4_sll_482_M1_6_115 ( .A(u4_sll_482_ML_int_6__115_), .B(
        u4_sll_482_ML_int_6__51_), .S(u4_sll_482_n42), .Z(
        u4_sll_482_ML_int_7__115_) );
  MUX2_X2 u4_sll_482_M1_6_116 ( .A(u4_sll_482_ML_int_6__116_), .B(
        u4_sll_482_ML_int_6__52_), .S(u4_sll_482_n42), .Z(
        u4_sll_482_ML_int_7__116_) );
  MUX2_X2 u4_sll_482_M1_6_117 ( .A(u4_sll_482_ML_int_6__117_), .B(
        u4_sll_482_ML_int_6__53_), .S(u4_sll_482_n42), .Z(
        u4_sll_482_ML_int_7__117_) );
  INV_X4 u4_sub_470_U27 ( .A(u4_fi_ldz_mi1_0_), .ZN(u4_sub_470_n16) );
  INV_X4 u4_sub_470_U26 ( .A(u4_fi_ldz_mi1_1_), .ZN(u4_sub_470_n15) );
  INV_X4 u4_sub_470_U25 ( .A(u4_fi_ldz_mi1_6_), .ZN(u4_sub_470_n14) );
  INV_X4 u4_sub_470_U24 ( .A(u4_fi_ldz_mi1_5_), .ZN(u4_sub_470_n13) );
  INV_X4 u4_sub_470_U23 ( .A(u4_fi_ldz_mi1_4_), .ZN(u4_sub_470_n12) );
  INV_X4 u4_sub_470_U22 ( .A(u4_fi_ldz_mi1_3_), .ZN(u4_sub_470_n11) );
  INV_X4 u4_sub_470_U21 ( .A(u4_fi_ldz_mi1_2_), .ZN(u4_sub_470_n10) );
  INV_X4 u4_sub_470_U20 ( .A(u4_exp_in_pl1_0_), .ZN(u4_sub_470_n9) );
  XNOR2_X2 u4_sub_470_U19 ( .A(u4_sub_470_n16), .B(u4_exp_in_pl1_0_), .ZN(
        u4_exp_next_mi_0_) );
  NAND2_X2 u4_sub_470_U18 ( .A1(u4_fi_ldz_mi1_0_), .A2(u4_sub_470_n9), .ZN(
        u4_sub_470_carry_1_) );
  INV_X4 u4_sub_470_U17 ( .A(u4_sub_470_carry_9_), .ZN(u4_sub_470_n8) );
  INV_X4 u4_sub_470_U16 ( .A(u4_exp_in_pl1_9_), .ZN(u4_sub_470_n7) );
  XNOR2_X2 u4_sub_470_U15 ( .A(u4_exp_in_pl1_9_), .B(u4_sub_470_carry_9_), 
        .ZN(u4_exp_next_mi_9_) );
  NAND2_X2 u4_sub_470_U14 ( .A1(u4_sub_470_n7), .A2(u4_sub_470_n8), .ZN(
        u4_sub_470_carry_10_) );
  INV_X4 u4_sub_470_U13 ( .A(u4_sub_470_carry_8_), .ZN(u4_sub_470_n6) );
  INV_X4 u4_sub_470_U12 ( .A(u4_exp_in_pl1_8_), .ZN(u4_sub_470_n5) );
  XNOR2_X2 u4_sub_470_U11 ( .A(u4_exp_in_pl1_8_), .B(u4_sub_470_carry_8_), 
        .ZN(u4_exp_next_mi_8_) );
  NAND2_X2 u4_sub_470_U10 ( .A1(u4_sub_470_n5), .A2(u4_sub_470_n6), .ZN(
        u4_sub_470_carry_9_) );
  INV_X4 u4_sub_470_U9 ( .A(u4_sub_470_carry_7_), .ZN(u4_sub_470_n4) );
  INV_X4 u4_sub_470_U8 ( .A(u4_exp_in_pl1_7_), .ZN(u4_sub_470_n3) );
  XNOR2_X2 u4_sub_470_U7 ( .A(u4_exp_in_pl1_7_), .B(u4_sub_470_carry_7_), .ZN(
        u4_exp_next_mi_7_) );
  NAND2_X2 u4_sub_470_U6 ( .A1(u4_sub_470_n3), .A2(u4_sub_470_n4), .ZN(
        u4_sub_470_carry_8_) );
  XNOR2_X2 u4_sub_470_U5 ( .A(u4_exp_in_pl1_11_), .B(u4_sub_470_carry_11_), 
        .ZN(u4_exp_next_mi_11_) );
  INV_X4 u4_sub_470_U4 ( .A(u4_sub_470_carry_10_), .ZN(u4_sub_470_n2) );
  INV_X4 u4_sub_470_U3 ( .A(u4_exp_in_pl1_10_), .ZN(u4_sub_470_n1) );
  XNOR2_X2 u4_sub_470_U2 ( .A(u4_exp_in_pl1_10_), .B(u4_sub_470_carry_10_), 
        .ZN(u4_exp_next_mi_10_) );
  NAND2_X2 u4_sub_470_U1 ( .A1(u4_sub_470_n1), .A2(u4_sub_470_n2), .ZN(
        u4_sub_470_carry_11_) );
  FA_X1 u4_sub_470_U2_1 ( .A(u4_exp_in_pl1_1_), .B(u4_sub_470_n15), .CI(
        u4_sub_470_carry_1_), .CO(u4_sub_470_carry_2_), .S(u4_exp_next_mi_1_)
         );
  FA_X1 u4_sub_470_U2_2 ( .A(u4_exp_in_pl1_2_), .B(u4_sub_470_n10), .CI(
        u4_sub_470_carry_2_), .CO(u4_sub_470_carry_3_), .S(u4_exp_next_mi_2_)
         );
  FA_X1 u4_sub_470_U2_3 ( .A(u4_exp_in_pl1_3_), .B(u4_sub_470_n11), .CI(
        u4_sub_470_carry_3_), .CO(u4_sub_470_carry_4_), .S(u4_exp_next_mi_3_)
         );
  FA_X1 u4_sub_470_U2_4 ( .A(u4_exp_in_pl1_4_), .B(u4_sub_470_n12), .CI(
        u4_sub_470_carry_4_), .CO(u4_sub_470_carry_5_), .S(u4_exp_next_mi_4_)
         );
  FA_X1 u4_sub_470_U2_5 ( .A(u4_exp_in_pl1_5_), .B(u4_sub_470_n13), .CI(
        u4_sub_470_carry_5_), .CO(u4_sub_470_carry_6_), .S(u4_exp_next_mi_5_)
         );
  FA_X1 u4_sub_470_U2_6 ( .A(u4_exp_in_pl1_6_), .B(u4_sub_470_n14), .CI(
        u4_sub_470_carry_6_), .CO(u4_sub_470_carry_7_), .S(u4_exp_next_mi_6_)
         );
  INV_X4 u4_sub_496_U23 ( .A(u4_ldz_all_0_), .ZN(u4_sub_496_n14) );
  INV_X4 u4_sub_496_U22 ( .A(u4_ldz_all_1_), .ZN(u4_sub_496_n13) );
  INV_X4 u4_sub_496_U21 ( .A(u4_ldz_all_2_), .ZN(u4_sub_496_n12) );
  INV_X4 u4_sub_496_U20 ( .A(u4_ldz_all_3_), .ZN(u4_sub_496_n11) );
  INV_X4 u4_sub_496_U19 ( .A(u4_ldz_all_4_), .ZN(u4_sub_496_n10) );
  INV_X4 u4_sub_496_U18 ( .A(u4_ldz_all_5_), .ZN(u4_sub_496_n9) );
  INV_X4 u4_sub_496_U17 ( .A(u4_ldz_all_6_), .ZN(u4_sub_496_n8) );
  INV_X4 u4_sub_496_U16 ( .A(u4_exp_in_pl1_0_), .ZN(u4_sub_496_n7) );
  XNOR2_X2 u4_sub_496_U15 ( .A(u4_sub_496_n14), .B(u4_exp_in_pl1_0_), .ZN(
        u4_div_exp2_0_) );
  NAND2_X2 u4_sub_496_U14 ( .A1(u4_ldz_all_0_), .A2(u4_sub_496_n7), .ZN(
        u4_sub_496_carry_1_) );
  INV_X4 u4_sub_496_U13 ( .A(u4_sub_496_carry_9_), .ZN(u4_sub_496_n6) );
  INV_X4 u4_sub_496_U12 ( .A(u4_exp_in_pl1_9_), .ZN(u4_sub_496_n5) );
  XNOR2_X2 u4_sub_496_U11 ( .A(u4_exp_in_pl1_9_), .B(u4_sub_496_carry_9_), 
        .ZN(u4_div_exp2_9_) );
  NAND2_X2 u4_sub_496_U10 ( .A1(u4_sub_496_n5), .A2(u4_sub_496_n6), .ZN(
        u4_sub_496_carry_10_) );
  INV_X4 u4_sub_496_U9 ( .A(u4_sub_496_carry_8_), .ZN(u4_sub_496_n4) );
  INV_X4 u4_sub_496_U8 ( .A(u4_exp_in_pl1_8_), .ZN(u4_sub_496_n3) );
  XNOR2_X2 u4_sub_496_U7 ( .A(u4_exp_in_pl1_8_), .B(u4_sub_496_carry_8_), .ZN(
        u4_div_exp2_8_) );
  NAND2_X2 u4_sub_496_U6 ( .A1(u4_sub_496_n3), .A2(u4_sub_496_n4), .ZN(
        u4_sub_496_carry_9_) );
  INV_X4 u4_sub_496_U5 ( .A(u4_sub_496_carry_7_), .ZN(u4_sub_496_n2) );
  INV_X4 u4_sub_496_U4 ( .A(u4_exp_in_pl1_7_), .ZN(u4_sub_496_n1) );
  XNOR2_X2 u4_sub_496_U3 ( .A(u4_exp_in_pl1_7_), .B(u4_sub_496_carry_7_), .ZN(
        u4_div_exp2_7_) );
  NAND2_X2 u4_sub_496_U2 ( .A1(u4_sub_496_n1), .A2(u4_sub_496_n2), .ZN(
        u4_sub_496_carry_8_) );
  XNOR2_X2 u4_sub_496_U1 ( .A(u4_exp_in_pl1_10_), .B(u4_sub_496_carry_10_), 
        .ZN(u4_div_exp2_10_) );
  FA_X1 u4_sub_496_U2_1 ( .A(u4_exp_in_pl1_1_), .B(u4_sub_496_n13), .CI(
        u4_sub_496_carry_1_), .CO(u4_sub_496_carry_2_), .S(u4_div_exp2_1_) );
  FA_X1 u4_sub_496_U2_2 ( .A(u4_exp_in_pl1_2_), .B(u4_sub_496_n12), .CI(
        u4_sub_496_carry_2_), .CO(u4_sub_496_carry_3_), .S(u4_div_exp2_2_) );
  FA_X1 u4_sub_496_U2_3 ( .A(u4_exp_in_pl1_3_), .B(u4_sub_496_n11), .CI(
        u4_sub_496_carry_3_), .CO(u4_sub_496_carry_4_), .S(u4_div_exp2_3_) );
  FA_X1 u4_sub_496_U2_4 ( .A(u4_exp_in_pl1_4_), .B(u4_sub_496_n10), .CI(
        u4_sub_496_carry_4_), .CO(u4_sub_496_carry_5_), .S(u4_div_exp2_4_) );
  FA_X1 u4_sub_496_U2_5 ( .A(u4_exp_in_pl1_5_), .B(u4_sub_496_n9), .CI(
        u4_sub_496_carry_5_), .CO(u4_sub_496_carry_6_), .S(u4_div_exp2_5_) );
  FA_X1 u4_sub_496_U2_6 ( .A(u4_exp_in_pl1_6_), .B(u4_sub_496_n8), .CI(
        u4_sub_496_carry_6_), .CO(u4_sub_496_carry_7_), .S(u4_div_exp2_6_) );
  AND2_X4 u4_add_489_U5 ( .A1(u4_fi_ldz_5_), .A2(u4_add_489_carry_5_), .ZN(
        u4_add_489_n5) );
  XOR2_X2 u4_add_489_U4 ( .A(u4_fi_ldz_5_), .B(u4_add_489_carry_5_), .Z(
        u4_ldz_all_5_) );
  AND2_X4 u4_add_489_U3 ( .A1(u4_fi_ldz_2a_0_), .A2(div_opa_ldz_r2[0]), .ZN(
        u4_add_489_n3) );
  XOR2_X2 u4_add_489_U2 ( .A(u4_fi_ldz_6_), .B(u4_add_489_n5), .Z(
        u4_ldz_all_6_) );
  XOR2_X2 u4_add_489_U1 ( .A(u4_fi_ldz_2a_0_), .B(div_opa_ldz_r2[0]), .Z(
        u4_ldz_all_0_) );
  FA_X1 u4_add_489_U1_1 ( .A(div_opa_ldz_r2[1]), .B(u4_fi_ldz_1_), .CI(
        u4_add_489_n3), .CO(u4_add_489_carry_2_), .S(u4_ldz_all_1_) );
  FA_X1 u4_add_489_U1_2 ( .A(div_opa_ldz_r2[2]), .B(u4_fi_ldz_2_), .CI(
        u4_add_489_carry_2_), .CO(u4_add_489_carry_3_), .S(u4_ldz_all_2_) );
  FA_X1 u4_add_489_U1_3 ( .A(div_opa_ldz_r2[3]), .B(u4_fi_ldz_3_), .CI(
        u4_add_489_carry_3_), .CO(u4_add_489_carry_4_), .S(u4_ldz_all_3_) );
  FA_X1 u4_add_489_U1_4 ( .A(div_opa_ldz_r2[4]), .B(u4_fi_ldz_4_), .CI(
        u4_add_489_carry_4_), .CO(u4_add_489_carry_5_), .S(u4_ldz_all_4_) );
  INV_X4 u4_add_466_U1 ( .A(n4600), .ZN(u4_exp_in_pl1_0_) );
  HA_X1 u4_add_466_U1_1_1 ( .A(exp_r[1]), .B(n4600), .CO(u4_add_466_carry[2]), 
        .S(u4_exp_in_pl1_1_) );
  HA_X1 u4_add_466_U1_1_2 ( .A(n4315), .B(u4_add_466_carry[2]), .CO(
        u4_add_466_carry[3]), .S(u4_exp_in_pl1_2_) );
  HA_X1 u4_add_466_U1_1_3 ( .A(n4655), .B(u4_add_466_carry[3]), .CO(
        u4_add_466_carry[4]), .S(u4_exp_in_pl1_3_) );
  HA_X1 u4_add_466_U1_1_4 ( .A(n4282), .B(u4_add_466_carry[4]), .CO(
        u4_add_466_carry[5]), .S(u4_exp_in_pl1_4_) );
  HA_X1 u4_add_466_U1_1_5 ( .A(n4290), .B(u4_add_466_carry[5]), .CO(
        u4_add_466_carry[6]), .S(u4_exp_in_pl1_5_) );
  HA_X1 u4_add_466_U1_1_6 ( .A(exp_r[6]), .B(u4_add_466_carry[6]), .CO(
        u4_add_466_carry[7]), .S(u4_exp_in_pl1_6_) );
  HA_X1 u4_add_466_U1_1_7 ( .A(n4281), .B(u4_add_466_carry[7]), .CO(
        u4_add_466_carry[8]), .S(u4_exp_in_pl1_7_) );
  HA_X1 u4_add_466_U1_1_8 ( .A(n4353), .B(u4_add_466_carry[8]), .CO(
        u4_add_466_carry[9]), .S(u4_exp_in_pl1_8_) );
  HA_X1 u4_add_466_U1_1_9 ( .A(n4289), .B(u4_add_466_carry[9]), .CO(
        u4_add_466_carry[10]), .S(u4_exp_in_pl1_9_) );
  HA_X1 u4_add_466_U1_1_10 ( .A(n4656), .B(u4_add_466_carry[10]), .CO(
        u4_exp_in_pl1_11_), .S(u4_exp_in_pl1_10_) );
  XOR2_X2 u4_add_494_U7 ( .A(u4_fi_ldz_2a_0_), .B(n4349), .Z(u4_div_exp1_0_)
         );
  AND2_X4 u4_add_494_U6 ( .A1(u4_exp_in_mi1_9_), .A2(u4_add_494_n5), .ZN(
        u4_add_494_n6) );
  AND2_X4 u4_add_494_U5 ( .A1(u4_exp_in_mi1_8_), .A2(u4_add_494_carry_8_), 
        .ZN(u4_add_494_n5) );
  AND2_X4 u4_add_494_U4 ( .A1(u4_fi_ldz_2a_0_), .A2(n4349), .ZN(u4_add_494_n4)
         );
  XOR2_X2 u4_add_494_U3 ( .A(u4_exp_in_mi1_8_), .B(u4_add_494_carry_8_), .Z(
        u4_div_exp1_8_) );
  XOR2_X2 u4_add_494_U2 ( .A(u4_exp_in_mi1_10_), .B(u4_add_494_n6), .Z(
        u4_div_exp1_10_) );
  XOR2_X2 u4_add_494_U1 ( .A(u4_exp_in_mi1_9_), .B(u4_add_494_n5), .Z(
        u4_div_exp1_9_) );
  FA_X1 u4_add_494_U1_1 ( .A(u4_exp_in_mi1_1_), .B(u4_fi_ldz_2a_1_), .CI(
        u4_add_494_n4), .CO(u4_add_494_carry_2_), .S(u4_div_exp1_1_) );
  FA_X1 u4_add_494_U1_2 ( .A(u4_exp_in_mi1_2_), .B(u4_fi_ldz_2a_2_), .CI(
        u4_add_494_carry_2_), .CO(u4_add_494_carry_3_), .S(u4_div_exp1_2_) );
  FA_X1 u4_add_494_U1_3 ( .A(u4_exp_in_mi1_3_), .B(u4_fi_ldz_2a_3_), .CI(
        u4_add_494_carry_3_), .CO(u4_add_494_carry_4_), .S(u4_div_exp1_3_) );
  FA_X1 u4_add_494_U1_4 ( .A(u4_exp_in_mi1_4_), .B(u4_fi_ldz_2a_4_), .CI(
        u4_add_494_carry_4_), .CO(u4_add_494_carry_5_), .S(u4_div_exp1_4_) );
  FA_X1 u4_add_494_U1_5 ( .A(u4_exp_in_mi1_5_), .B(u4_fi_ldz_2a_5_), .CI(
        u4_add_494_carry_5_), .CO(u4_add_494_carry_6_), .S(u4_div_exp1_5_) );
  FA_X1 u4_add_494_U1_6 ( .A(u4_exp_in_mi1_6_), .B(u4_fi_ldz_2a_6_), .CI(
        u4_add_494_carry_6_), .CO(u4_add_494_carry_7_), .S(u4_div_exp1_6_) );
  FA_X1 u4_add_494_U1_7 ( .A(u4_exp_in_mi1_7_), .B(u4_fi_ldz_2a_6_), .CI(
        u4_add_494_carry_7_), .CO(u4_add_494_carry_8_), .S(u4_div_exp1_7_) );
  INV_X1 u4_add_396_U1 ( .A(u4_fract_out_0_), .ZN(u4_fract_out_pl1_0_) );
  HA_X1 u4_add_396_U1_1_1 ( .A(u4_fract_out_1_), .B(u4_fract_out_0_), .CO(
        u4_add_396_carry[2]), .S(u4_fract_out_pl1_1_) );
  HA_X1 u4_add_396_U1_1_2 ( .A(u4_fract_out_2_), .B(u4_add_396_carry[2]), .CO(
        u4_add_396_carry[3]), .S(u4_fract_out_pl1_2_) );
  HA_X1 u4_add_396_U1_1_3 ( .A(u4_fract_out_3_), .B(u4_add_396_carry[3]), .CO(
        u4_add_396_carry[4]), .S(u4_fract_out_pl1_3_) );
  HA_X1 u4_add_396_U1_1_4 ( .A(u4_fract_out_4_), .B(u4_add_396_carry[4]), .CO(
        u4_add_396_carry[5]), .S(u4_fract_out_pl1_4_) );
  HA_X1 u4_add_396_U1_1_5 ( .A(u4_fract_out_5_), .B(u4_add_396_carry[5]), .CO(
        u4_add_396_carry[6]), .S(u4_fract_out_pl1_5_) );
  HA_X1 u4_add_396_U1_1_6 ( .A(u4_fract_out_6_), .B(u4_add_396_carry[6]), .CO(
        u4_add_396_carry[7]), .S(u4_fract_out_pl1_6_) );
  HA_X1 u4_add_396_U1_1_7 ( .A(u4_fract_out_7_), .B(u4_add_396_carry[7]), .CO(
        u4_add_396_carry[8]), .S(u4_fract_out_pl1_7_) );
  HA_X1 u4_add_396_U1_1_8 ( .A(u4_fract_out_8_), .B(u4_add_396_carry[8]), .CO(
        u4_add_396_carry[9]), .S(u4_fract_out_pl1_8_) );
  HA_X1 u4_add_396_U1_1_9 ( .A(u4_fract_out_9_), .B(u4_add_396_carry[9]), .CO(
        u4_add_396_carry[10]), .S(u4_fract_out_pl1_9_) );
  HA_X1 u4_add_396_U1_1_10 ( .A(u4_fract_out_10_), .B(u4_add_396_carry[10]), 
        .CO(u4_add_396_carry[11]), .S(u4_fract_out_pl1_10_) );
  HA_X1 u4_add_396_U1_1_11 ( .A(u4_fract_out_11_), .B(u4_add_396_carry[11]), 
        .CO(u4_add_396_carry[12]), .S(u4_fract_out_pl1_11_) );
  HA_X1 u4_add_396_U1_1_12 ( .A(u4_fract_out_12_), .B(u4_add_396_carry[12]), 
        .CO(u4_add_396_carry[13]), .S(u4_fract_out_pl1_12_) );
  HA_X1 u4_add_396_U1_1_13 ( .A(u4_fract_out_13_), .B(u4_add_396_carry[13]), 
        .CO(u4_add_396_carry[14]), .S(u4_fract_out_pl1_13_) );
  HA_X1 u4_add_396_U1_1_14 ( .A(u4_fract_out_14_), .B(u4_add_396_carry[14]), 
        .CO(u4_add_396_carry[15]), .S(u4_fract_out_pl1_14_) );
  HA_X1 u4_add_396_U1_1_15 ( .A(u4_fract_out_15_), .B(u4_add_396_carry[15]), 
        .CO(u4_add_396_carry[16]), .S(u4_fract_out_pl1_15_) );
  HA_X1 u4_add_396_U1_1_16 ( .A(u4_fract_out_16_), .B(u4_add_396_carry[16]), 
        .CO(u4_add_396_carry[17]), .S(u4_fract_out_pl1_16_) );
  HA_X1 u4_add_396_U1_1_17 ( .A(u4_fract_out_17_), .B(u4_add_396_carry[17]), 
        .CO(u4_add_396_carry[18]), .S(u4_fract_out_pl1_17_) );
  HA_X1 u4_add_396_U1_1_18 ( .A(u4_fract_out_18_), .B(u4_add_396_carry[18]), 
        .CO(u4_add_396_carry[19]), .S(u4_fract_out_pl1_18_) );
  HA_X1 u4_add_396_U1_1_19 ( .A(u4_fract_out_19_), .B(u4_add_396_carry[19]), 
        .CO(u4_add_396_carry[20]), .S(u4_fract_out_pl1_19_) );
  HA_X1 u4_add_396_U1_1_20 ( .A(u4_fract_out_20_), .B(u4_add_396_carry[20]), 
        .CO(u4_add_396_carry[21]), .S(u4_fract_out_pl1_20_) );
  HA_X1 u4_add_396_U1_1_21 ( .A(u4_fract_out_21_), .B(u4_add_396_carry[21]), 
        .CO(u4_add_396_carry[22]), .S(u4_fract_out_pl1_21_) );
  HA_X1 u4_add_396_U1_1_22 ( .A(u4_fract_out_22_), .B(u4_add_396_carry[22]), 
        .CO(u4_add_396_carry[23]), .S(u4_fract_out_pl1_22_) );
  HA_X1 u4_add_396_U1_1_23 ( .A(u4_fract_out_23_), .B(u4_add_396_carry[23]), 
        .CO(u4_add_396_carry[24]), .S(u4_fract_out_pl1_23_) );
  HA_X1 u4_add_396_U1_1_24 ( .A(u4_fract_out_24_), .B(u4_add_396_carry[24]), 
        .CO(u4_add_396_carry[25]), .S(u4_fract_out_pl1_24_) );
  HA_X1 u4_add_396_U1_1_25 ( .A(u4_fract_out_25_), .B(u4_add_396_carry[25]), 
        .CO(u4_add_396_carry[26]), .S(u4_fract_out_pl1_25_) );
  HA_X1 u4_add_396_U1_1_26 ( .A(u4_fract_out_26_), .B(u4_add_396_carry[26]), 
        .CO(u4_add_396_carry[27]), .S(u4_fract_out_pl1_26_) );
  HA_X1 u4_add_396_U1_1_27 ( .A(u4_fract_out_27_), .B(u4_add_396_carry[27]), 
        .CO(u4_add_396_carry[28]), .S(u4_fract_out_pl1_27_) );
  HA_X1 u4_add_396_U1_1_28 ( .A(u4_fract_out_28_), .B(u4_add_396_carry[28]), 
        .CO(u4_add_396_carry[29]), .S(u4_fract_out_pl1_28_) );
  HA_X1 u4_add_396_U1_1_29 ( .A(u4_fract_out_29_), .B(u4_add_396_carry[29]), 
        .CO(u4_add_396_carry[30]), .S(u4_fract_out_pl1_29_) );
  HA_X1 u4_add_396_U1_1_30 ( .A(u4_fract_out_30_), .B(u4_add_396_carry[30]), 
        .CO(u4_add_396_carry[31]), .S(u4_fract_out_pl1_30_) );
  HA_X1 u4_add_396_U1_1_31 ( .A(u4_fract_out_31_), .B(u4_add_396_carry[31]), 
        .CO(u4_add_396_carry[32]), .S(u4_fract_out_pl1_31_) );
  HA_X1 u4_add_396_U1_1_32 ( .A(u4_fract_out_32_), .B(u4_add_396_carry[32]), 
        .CO(u4_add_396_carry[33]), .S(u4_fract_out_pl1_32_) );
  HA_X1 u4_add_396_U1_1_33 ( .A(u4_fract_out_33_), .B(u4_add_396_carry[33]), 
        .CO(u4_add_396_carry[34]), .S(u4_fract_out_pl1_33_) );
  HA_X1 u4_add_396_U1_1_34 ( .A(u4_fract_out_34_), .B(u4_add_396_carry[34]), 
        .CO(u4_add_396_carry[35]), .S(u4_fract_out_pl1_34_) );
  HA_X1 u4_add_396_U1_1_35 ( .A(u4_fract_out_35_), .B(u4_add_396_carry[35]), 
        .CO(u4_add_396_carry[36]), .S(u4_fract_out_pl1_35_) );
  HA_X1 u4_add_396_U1_1_36 ( .A(u4_fract_out_36_), .B(u4_add_396_carry[36]), 
        .CO(u4_add_396_carry[37]), .S(u4_fract_out_pl1_36_) );
  HA_X1 u4_add_396_U1_1_37 ( .A(u4_fract_out_37_), .B(u4_add_396_carry[37]), 
        .CO(u4_add_396_carry[38]), .S(u4_fract_out_pl1_37_) );
  HA_X1 u4_add_396_U1_1_38 ( .A(u4_fract_out_38_), .B(u4_add_396_carry[38]), 
        .CO(u4_add_396_carry[39]), .S(u4_fract_out_pl1_38_) );
  HA_X1 u4_add_396_U1_1_39 ( .A(u4_fract_out_39_), .B(u4_add_396_carry[39]), 
        .CO(u4_add_396_carry[40]), .S(u4_fract_out_pl1_39_) );
  HA_X1 u4_add_396_U1_1_40 ( .A(u4_fract_out_40_), .B(u4_add_396_carry[40]), 
        .CO(u4_add_396_carry[41]), .S(u4_fract_out_pl1_40_) );
  HA_X1 u4_add_396_U1_1_41 ( .A(u4_fract_out_41_), .B(u4_add_396_carry[41]), 
        .CO(u4_add_396_carry[42]), .S(u4_fract_out_pl1_41_) );
  HA_X1 u4_add_396_U1_1_42 ( .A(u4_fract_out_42_), .B(u4_add_396_carry[42]), 
        .CO(u4_add_396_carry[43]), .S(u4_fract_out_pl1_42_) );
  HA_X1 u4_add_396_U1_1_43 ( .A(u4_fract_out_43_), .B(u4_add_396_carry[43]), 
        .CO(u4_add_396_carry[44]), .S(u4_fract_out_pl1_43_) );
  HA_X1 u4_add_396_U1_1_44 ( .A(u4_fract_out_44_), .B(u4_add_396_carry[44]), 
        .CO(u4_add_396_carry[45]), .S(u4_fract_out_pl1_44_) );
  HA_X1 u4_add_396_U1_1_45 ( .A(u4_fract_out_45_), .B(u4_add_396_carry[45]), 
        .CO(u4_add_396_carry[46]), .S(u4_fract_out_pl1_45_) );
  HA_X1 u4_add_396_U1_1_46 ( .A(u4_fract_out_46_), .B(u4_add_396_carry[46]), 
        .CO(u4_add_396_carry[47]), .S(u4_fract_out_pl1_46_) );
  HA_X1 u4_add_396_U1_1_47 ( .A(u4_fract_out_47_), .B(u4_add_396_carry[47]), 
        .CO(u4_add_396_carry[48]), .S(u4_fract_out_pl1_47_) );
  HA_X1 u4_add_396_U1_1_48 ( .A(u4_fract_out_48_), .B(u4_add_396_carry[48]), 
        .CO(u4_add_396_carry[49]), .S(u4_fract_out_pl1_48_) );
  HA_X1 u4_add_396_U1_1_49 ( .A(u4_fract_out_49_), .B(u4_add_396_carry[49]), 
        .CO(u4_add_396_carry[50]), .S(u4_fract_out_pl1_49_) );
  HA_X1 u4_add_396_U1_1_50 ( .A(u4_fract_out_50_), .B(u4_add_396_carry[50]), 
        .CO(u4_add_396_carry[51]), .S(u4_fract_out_pl1_50_) );
  HA_X1 u4_add_396_U1_1_51 ( .A(u4_fract_out_51_), .B(u4_add_396_carry[51]), 
        .CO(u4_fract_out_pl1_52_), .S(u4_fract_out_pl1_51_) );
  INV_X4 u3_sub_63_U60 ( .A(fractb[55]), .ZN(u3_sub_63_n58) );
  INV_X4 u3_sub_63_U59 ( .A(fractb[54]), .ZN(u3_sub_63_n57) );
  INV_X4 u3_sub_63_U58 ( .A(fractb[53]), .ZN(u3_sub_63_n56) );
  INV_X4 u3_sub_63_U57 ( .A(fractb[52]), .ZN(u3_sub_63_n55) );
  INV_X4 u3_sub_63_U56 ( .A(fractb[51]), .ZN(u3_sub_63_n54) );
  INV_X4 u3_sub_63_U55 ( .A(fractb[50]), .ZN(u3_sub_63_n53) );
  INV_X4 u3_sub_63_U54 ( .A(fractb[49]), .ZN(u3_sub_63_n52) );
  INV_X4 u3_sub_63_U53 ( .A(fractb[48]), .ZN(u3_sub_63_n51) );
  INV_X4 u3_sub_63_U52 ( .A(fractb[47]), .ZN(u3_sub_63_n50) );
  INV_X4 u3_sub_63_U51 ( .A(fractb[46]), .ZN(u3_sub_63_n49) );
  INV_X4 u3_sub_63_U50 ( .A(fractb[45]), .ZN(u3_sub_63_n48) );
  INV_X4 u3_sub_63_U49 ( .A(fractb[44]), .ZN(u3_sub_63_n47) );
  INV_X4 u3_sub_63_U48 ( .A(fractb[43]), .ZN(u3_sub_63_n46) );
  INV_X4 u3_sub_63_U47 ( .A(fractb[42]), .ZN(u3_sub_63_n45) );
  INV_X4 u3_sub_63_U46 ( .A(fractb[41]), .ZN(u3_sub_63_n44) );
  INV_X4 u3_sub_63_U45 ( .A(fractb[40]), .ZN(u3_sub_63_n43) );
  INV_X4 u3_sub_63_U44 ( .A(fractb[39]), .ZN(u3_sub_63_n42) );
  INV_X4 u3_sub_63_U43 ( .A(fractb[38]), .ZN(u3_sub_63_n41) );
  INV_X4 u3_sub_63_U42 ( .A(fractb[37]), .ZN(u3_sub_63_n40) );
  INV_X4 u3_sub_63_U41 ( .A(fractb[36]), .ZN(u3_sub_63_n39) );
  INV_X4 u3_sub_63_U40 ( .A(fractb[35]), .ZN(u3_sub_63_n38) );
  INV_X4 u3_sub_63_U39 ( .A(fractb[34]), .ZN(u3_sub_63_n37) );
  INV_X4 u3_sub_63_U38 ( .A(fractb[33]), .ZN(u3_sub_63_n36) );
  INV_X4 u3_sub_63_U37 ( .A(fractb[32]), .ZN(u3_sub_63_n35) );
  INV_X4 u3_sub_63_U36 ( .A(fractb[31]), .ZN(u3_sub_63_n34) );
  INV_X4 u3_sub_63_U35 ( .A(fractb[30]), .ZN(u3_sub_63_n33) );
  INV_X4 u3_sub_63_U34 ( .A(fractb[29]), .ZN(u3_sub_63_n32) );
  INV_X4 u3_sub_63_U33 ( .A(fractb[28]), .ZN(u3_sub_63_n31) );
  INV_X4 u3_sub_63_U32 ( .A(fractb[27]), .ZN(u3_sub_63_n30) );
  INV_X4 u3_sub_63_U31 ( .A(fractb[26]), .ZN(u3_sub_63_n29) );
  INV_X4 u3_sub_63_U30 ( .A(fractb[25]), .ZN(u3_sub_63_n28) );
  INV_X4 u3_sub_63_U29 ( .A(fractb[24]), .ZN(u3_sub_63_n27) );
  INV_X4 u3_sub_63_U28 ( .A(fractb[23]), .ZN(u3_sub_63_n26) );
  INV_X4 u3_sub_63_U27 ( .A(fractb[22]), .ZN(u3_sub_63_n25) );
  INV_X4 u3_sub_63_U26 ( .A(fractb[21]), .ZN(u3_sub_63_n24) );
  INV_X4 u3_sub_63_U25 ( .A(fractb[20]), .ZN(u3_sub_63_n23) );
  INV_X4 u3_sub_63_U24 ( .A(fractb[19]), .ZN(u3_sub_63_n22) );
  INV_X4 u3_sub_63_U23 ( .A(fractb[18]), .ZN(u3_sub_63_n21) );
  INV_X4 u3_sub_63_U22 ( .A(fractb[17]), .ZN(u3_sub_63_n20) );
  INV_X4 u3_sub_63_U21 ( .A(fractb[16]), .ZN(u3_sub_63_n19) );
  INV_X4 u3_sub_63_U20 ( .A(fractb[15]), .ZN(u3_sub_63_n18) );
  INV_X4 u3_sub_63_U19 ( .A(fractb[14]), .ZN(u3_sub_63_n17) );
  INV_X4 u3_sub_63_U18 ( .A(fractb[13]), .ZN(u3_sub_63_n16) );
  INV_X4 u3_sub_63_U17 ( .A(fractb[12]), .ZN(u3_sub_63_n15) );
  INV_X4 u3_sub_63_U16 ( .A(fractb[11]), .ZN(u3_sub_63_n14) );
  INV_X4 u3_sub_63_U15 ( .A(fractb[10]), .ZN(u3_sub_63_n13) );
  INV_X4 u3_sub_63_U14 ( .A(fractb[9]), .ZN(u3_sub_63_n12) );
  INV_X4 u3_sub_63_U13 ( .A(fractb[8]), .ZN(u3_sub_63_n11) );
  INV_X4 u3_sub_63_U12 ( .A(fractb[7]), .ZN(u3_sub_63_n10) );
  INV_X4 u3_sub_63_U11 ( .A(fractb[6]), .ZN(u3_sub_63_n9) );
  INV_X4 u3_sub_63_U10 ( .A(fractb[5]), .ZN(u3_sub_63_n8) );
  INV_X4 u3_sub_63_U9 ( .A(fractb[4]), .ZN(u3_sub_63_n7) );
  INV_X4 u3_sub_63_U8 ( .A(fractb[3]), .ZN(u3_sub_63_n6) );
  INV_X4 u3_sub_63_U7 ( .A(fractb[2]), .ZN(u3_sub_63_n5) );
  INV_X4 u3_sub_63_U6 ( .A(fractb[1]), .ZN(u3_sub_63_n4) );
  INV_X4 u3_sub_63_U5 ( .A(fractb[0]), .ZN(u3_sub_63_n3) );
  INV_X4 u3_sub_63_U4 ( .A(u3_sub_63_carry[56]), .ZN(u3_N116) );
  INV_X4 u3_sub_63_U3 ( .A(fracta[0]), .ZN(u3_sub_63_n1) );
  XNOR2_X2 u3_sub_63_U2 ( .A(u3_sub_63_n3), .B(fracta[0]), .ZN(u3_N60) );
  NAND2_X2 u3_sub_63_U1 ( .A1(fractb[0]), .A2(u3_sub_63_n1), .ZN(
        u3_sub_63_carry[1]) );
  FA_X1 u3_sub_63_U2_1 ( .A(fracta[1]), .B(u3_sub_63_n4), .CI(
        u3_sub_63_carry[1]), .CO(u3_sub_63_carry[2]), .S(u3_N61) );
  FA_X1 u3_sub_63_U2_2 ( .A(fracta[2]), .B(u3_sub_63_n5), .CI(
        u3_sub_63_carry[2]), .CO(u3_sub_63_carry[3]), .S(u3_N62) );
  FA_X1 u3_sub_63_U2_3 ( .A(fracta[3]), .B(u3_sub_63_n6), .CI(
        u3_sub_63_carry[3]), .CO(u3_sub_63_carry[4]), .S(u3_N63) );
  FA_X1 u3_sub_63_U2_4 ( .A(fracta[4]), .B(u3_sub_63_n7), .CI(
        u3_sub_63_carry[4]), .CO(u3_sub_63_carry[5]), .S(u3_N64) );
  FA_X1 u3_sub_63_U2_5 ( .A(fracta[5]), .B(u3_sub_63_n8), .CI(
        u3_sub_63_carry[5]), .CO(u3_sub_63_carry[6]), .S(u3_N65) );
  FA_X1 u3_sub_63_U2_6 ( .A(fracta[6]), .B(u3_sub_63_n9), .CI(
        u3_sub_63_carry[6]), .CO(u3_sub_63_carry[7]), .S(u3_N66) );
  FA_X1 u3_sub_63_U2_7 ( .A(fracta[7]), .B(u3_sub_63_n10), .CI(
        u3_sub_63_carry[7]), .CO(u3_sub_63_carry[8]), .S(u3_N67) );
  FA_X1 u3_sub_63_U2_8 ( .A(fracta[8]), .B(u3_sub_63_n11), .CI(
        u3_sub_63_carry[8]), .CO(u3_sub_63_carry[9]), .S(u3_N68) );
  FA_X1 u3_sub_63_U2_9 ( .A(fracta[9]), .B(u3_sub_63_n12), .CI(
        u3_sub_63_carry[9]), .CO(u3_sub_63_carry[10]), .S(u3_N69) );
  FA_X1 u3_sub_63_U2_10 ( .A(fracta[10]), .B(u3_sub_63_n13), .CI(
        u3_sub_63_carry[10]), .CO(u3_sub_63_carry[11]), .S(u3_N70) );
  FA_X1 u3_sub_63_U2_11 ( .A(fracta[11]), .B(u3_sub_63_n14), .CI(
        u3_sub_63_carry[11]), .CO(u3_sub_63_carry[12]), .S(u3_N71) );
  FA_X1 u3_sub_63_U2_12 ( .A(fracta[12]), .B(u3_sub_63_n15), .CI(
        u3_sub_63_carry[12]), .CO(u3_sub_63_carry[13]), .S(u3_N72) );
  FA_X1 u3_sub_63_U2_13 ( .A(fracta[13]), .B(u3_sub_63_n16), .CI(
        u3_sub_63_carry[13]), .CO(u3_sub_63_carry[14]), .S(u3_N73) );
  FA_X1 u3_sub_63_U2_14 ( .A(fracta[14]), .B(u3_sub_63_n17), .CI(
        u3_sub_63_carry[14]), .CO(u3_sub_63_carry[15]), .S(u3_N74) );
  FA_X1 u3_sub_63_U2_15 ( .A(fracta[15]), .B(u3_sub_63_n18), .CI(
        u3_sub_63_carry[15]), .CO(u3_sub_63_carry[16]), .S(u3_N75) );
  FA_X1 u3_sub_63_U2_16 ( .A(fracta[16]), .B(u3_sub_63_n19), .CI(
        u3_sub_63_carry[16]), .CO(u3_sub_63_carry[17]), .S(u3_N76) );
  FA_X1 u3_sub_63_U2_17 ( .A(fracta[17]), .B(u3_sub_63_n20), .CI(
        u3_sub_63_carry[17]), .CO(u3_sub_63_carry[18]), .S(u3_N77) );
  FA_X1 u3_sub_63_U2_18 ( .A(fracta[18]), .B(u3_sub_63_n21), .CI(
        u3_sub_63_carry[18]), .CO(u3_sub_63_carry[19]), .S(u3_N78) );
  FA_X1 u3_sub_63_U2_19 ( .A(fracta[19]), .B(u3_sub_63_n22), .CI(
        u3_sub_63_carry[19]), .CO(u3_sub_63_carry[20]), .S(u3_N79) );
  FA_X1 u3_sub_63_U2_20 ( .A(fracta[20]), .B(u3_sub_63_n23), .CI(
        u3_sub_63_carry[20]), .CO(u3_sub_63_carry[21]), .S(u3_N80) );
  FA_X1 u3_sub_63_U2_21 ( .A(fracta[21]), .B(u3_sub_63_n24), .CI(
        u3_sub_63_carry[21]), .CO(u3_sub_63_carry[22]), .S(u3_N81) );
  FA_X1 u3_sub_63_U2_22 ( .A(fracta[22]), .B(u3_sub_63_n25), .CI(
        u3_sub_63_carry[22]), .CO(u3_sub_63_carry[23]), .S(u3_N82) );
  FA_X1 u3_sub_63_U2_23 ( .A(fracta[23]), .B(u3_sub_63_n26), .CI(
        u3_sub_63_carry[23]), .CO(u3_sub_63_carry[24]), .S(u3_N83) );
  FA_X1 u3_sub_63_U2_24 ( .A(fracta[24]), .B(u3_sub_63_n27), .CI(
        u3_sub_63_carry[24]), .CO(u3_sub_63_carry[25]), .S(u3_N84) );
  FA_X1 u3_sub_63_U2_25 ( .A(fracta[25]), .B(u3_sub_63_n28), .CI(
        u3_sub_63_carry[25]), .CO(u3_sub_63_carry[26]), .S(u3_N85) );
  FA_X1 u3_sub_63_U2_26 ( .A(fracta[26]), .B(u3_sub_63_n29), .CI(
        u3_sub_63_carry[26]), .CO(u3_sub_63_carry[27]), .S(u3_N86) );
  FA_X1 u3_sub_63_U2_27 ( .A(fracta[27]), .B(u3_sub_63_n30), .CI(
        u3_sub_63_carry[27]), .CO(u3_sub_63_carry[28]), .S(u3_N87) );
  FA_X1 u3_sub_63_U2_28 ( .A(fracta[28]), .B(u3_sub_63_n31), .CI(
        u3_sub_63_carry[28]), .CO(u3_sub_63_carry[29]), .S(u3_N88) );
  FA_X1 u3_sub_63_U2_29 ( .A(fracta[29]), .B(u3_sub_63_n32), .CI(
        u3_sub_63_carry[29]), .CO(u3_sub_63_carry[30]), .S(u3_N89) );
  FA_X1 u3_sub_63_U2_30 ( .A(fracta[30]), .B(u3_sub_63_n33), .CI(
        u3_sub_63_carry[30]), .CO(u3_sub_63_carry[31]), .S(u3_N90) );
  FA_X1 u3_sub_63_U2_31 ( .A(fracta[31]), .B(u3_sub_63_n34), .CI(
        u3_sub_63_carry[31]), .CO(u3_sub_63_carry[32]), .S(u3_N91) );
  FA_X1 u3_sub_63_U2_32 ( .A(fracta[32]), .B(u3_sub_63_n35), .CI(
        u3_sub_63_carry[32]), .CO(u3_sub_63_carry[33]), .S(u3_N92) );
  FA_X1 u3_sub_63_U2_33 ( .A(fracta[33]), .B(u3_sub_63_n36), .CI(
        u3_sub_63_carry[33]), .CO(u3_sub_63_carry[34]), .S(u3_N93) );
  FA_X1 u3_sub_63_U2_34 ( .A(fracta[34]), .B(u3_sub_63_n37), .CI(
        u3_sub_63_carry[34]), .CO(u3_sub_63_carry[35]), .S(u3_N94) );
  FA_X1 u3_sub_63_U2_35 ( .A(fracta[35]), .B(u3_sub_63_n38), .CI(
        u3_sub_63_carry[35]), .CO(u3_sub_63_carry[36]), .S(u3_N95) );
  FA_X1 u3_sub_63_U2_36 ( .A(fracta[36]), .B(u3_sub_63_n39), .CI(
        u3_sub_63_carry[36]), .CO(u3_sub_63_carry[37]), .S(u3_N96) );
  FA_X1 u3_sub_63_U2_37 ( .A(fracta[37]), .B(u3_sub_63_n40), .CI(
        u3_sub_63_carry[37]), .CO(u3_sub_63_carry[38]), .S(u3_N97) );
  FA_X1 u3_sub_63_U2_38 ( .A(fracta[38]), .B(u3_sub_63_n41), .CI(
        u3_sub_63_carry[38]), .CO(u3_sub_63_carry[39]), .S(u3_N98) );
  FA_X1 u3_sub_63_U2_39 ( .A(fracta[39]), .B(u3_sub_63_n42), .CI(
        u3_sub_63_carry[39]), .CO(u3_sub_63_carry[40]), .S(u3_N99) );
  FA_X1 u3_sub_63_U2_40 ( .A(fracta[40]), .B(u3_sub_63_n43), .CI(
        u3_sub_63_carry[40]), .CO(u3_sub_63_carry[41]), .S(u3_N100) );
  FA_X1 u3_sub_63_U2_41 ( .A(fracta[41]), .B(u3_sub_63_n44), .CI(
        u3_sub_63_carry[41]), .CO(u3_sub_63_carry[42]), .S(u3_N101) );
  FA_X1 u3_sub_63_U2_42 ( .A(fracta[42]), .B(u3_sub_63_n45), .CI(
        u3_sub_63_carry[42]), .CO(u3_sub_63_carry[43]), .S(u3_N102) );
  FA_X1 u3_sub_63_U2_43 ( .A(fracta[43]), .B(u3_sub_63_n46), .CI(
        u3_sub_63_carry[43]), .CO(u3_sub_63_carry[44]), .S(u3_N103) );
  FA_X1 u3_sub_63_U2_44 ( .A(fracta[44]), .B(u3_sub_63_n47), .CI(
        u3_sub_63_carry[44]), .CO(u3_sub_63_carry[45]), .S(u3_N104) );
  FA_X1 u3_sub_63_U2_45 ( .A(fracta[45]), .B(u3_sub_63_n48), .CI(
        u3_sub_63_carry[45]), .CO(u3_sub_63_carry[46]), .S(u3_N105) );
  FA_X1 u3_sub_63_U2_46 ( .A(fracta[46]), .B(u3_sub_63_n49), .CI(
        u3_sub_63_carry[46]), .CO(u3_sub_63_carry[47]), .S(u3_N106) );
  FA_X1 u3_sub_63_U2_47 ( .A(fracta[47]), .B(u3_sub_63_n50), .CI(
        u3_sub_63_carry[47]), .CO(u3_sub_63_carry[48]), .S(u3_N107) );
  FA_X1 u3_sub_63_U2_48 ( .A(fracta[48]), .B(u3_sub_63_n51), .CI(
        u3_sub_63_carry[48]), .CO(u3_sub_63_carry[49]), .S(u3_N108) );
  FA_X1 u3_sub_63_U2_49 ( .A(fracta[49]), .B(u3_sub_63_n52), .CI(
        u3_sub_63_carry[49]), .CO(u3_sub_63_carry[50]), .S(u3_N109) );
  FA_X1 u3_sub_63_U2_50 ( .A(fracta[50]), .B(u3_sub_63_n53), .CI(
        u3_sub_63_carry[50]), .CO(u3_sub_63_carry[51]), .S(u3_N110) );
  FA_X1 u3_sub_63_U2_51 ( .A(fracta[51]), .B(u3_sub_63_n54), .CI(
        u3_sub_63_carry[51]), .CO(u3_sub_63_carry[52]), .S(u3_N111) );
  FA_X1 u3_sub_63_U2_52 ( .A(fracta[52]), .B(u3_sub_63_n55), .CI(
        u3_sub_63_carry[52]), .CO(u3_sub_63_carry[53]), .S(u3_N112) );
  FA_X1 u3_sub_63_U2_53 ( .A(fracta[53]), .B(u3_sub_63_n56), .CI(
        u3_sub_63_carry[53]), .CO(u3_sub_63_carry[54]), .S(u3_N113) );
  FA_X1 u3_sub_63_U2_54 ( .A(fracta[54]), .B(u3_sub_63_n57), .CI(
        u3_sub_63_carry[54]), .CO(u3_sub_63_carry[55]), .S(u3_N114) );
  FA_X1 u3_sub_63_U2_55 ( .A(fracta[55]), .B(u3_sub_63_n58), .CI(
        u3_sub_63_carry[55]), .CO(u3_sub_63_carry[56]), .S(u3_N115) );
  AND2_X4 u3_add_63_U2 ( .A1(fractb[0]), .A2(fracta[0]), .ZN(u3_add_63_n2) );
  XOR2_X2 u3_add_63_U1 ( .A(fractb[0]), .B(fracta[0]), .Z(u3_N3) );
  FA_X1 u3_add_63_U1_1 ( .A(fracta[1]), .B(fractb[1]), .CI(u3_add_63_n2), .CO(
        u3_add_63_carry[2]), .S(u3_N4) );
  FA_X1 u3_add_63_U1_2 ( .A(fracta[2]), .B(fractb[2]), .CI(u3_add_63_carry[2]), 
        .CO(u3_add_63_carry[3]), .S(u3_N5) );
  FA_X1 u3_add_63_U1_3 ( .A(fracta[3]), .B(fractb[3]), .CI(u3_add_63_carry[3]), 
        .CO(u3_add_63_carry[4]), .S(u3_N6) );
  FA_X1 u3_add_63_U1_4 ( .A(fracta[4]), .B(fractb[4]), .CI(u3_add_63_carry[4]), 
        .CO(u3_add_63_carry[5]), .S(u3_N7) );
  FA_X1 u3_add_63_U1_5 ( .A(fracta[5]), .B(fractb[5]), .CI(u3_add_63_carry[5]), 
        .CO(u3_add_63_carry[6]), .S(u3_N8) );
  FA_X1 u3_add_63_U1_6 ( .A(fracta[6]), .B(fractb[6]), .CI(u3_add_63_carry[6]), 
        .CO(u3_add_63_carry[7]), .S(u3_N9) );
  FA_X1 u3_add_63_U1_7 ( .A(fracta[7]), .B(fractb[7]), .CI(u3_add_63_carry[7]), 
        .CO(u3_add_63_carry[8]), .S(u3_N10) );
  FA_X1 u3_add_63_U1_8 ( .A(fracta[8]), .B(fractb[8]), .CI(u3_add_63_carry[8]), 
        .CO(u3_add_63_carry[9]), .S(u3_N11) );
  FA_X1 u3_add_63_U1_9 ( .A(fracta[9]), .B(fractb[9]), .CI(u3_add_63_carry[9]), 
        .CO(u3_add_63_carry[10]), .S(u3_N12) );
  FA_X1 u3_add_63_U1_10 ( .A(fracta[10]), .B(fractb[10]), .CI(
        u3_add_63_carry[10]), .CO(u3_add_63_carry[11]), .S(u3_N13) );
  FA_X1 u3_add_63_U1_11 ( .A(fracta[11]), .B(fractb[11]), .CI(
        u3_add_63_carry[11]), .CO(u3_add_63_carry[12]), .S(u3_N14) );
  FA_X1 u3_add_63_U1_12 ( .A(fracta[12]), .B(fractb[12]), .CI(
        u3_add_63_carry[12]), .CO(u3_add_63_carry[13]), .S(u3_N15) );
  FA_X1 u3_add_63_U1_13 ( .A(fracta[13]), .B(fractb[13]), .CI(
        u3_add_63_carry[13]), .CO(u3_add_63_carry[14]), .S(u3_N16) );
  FA_X1 u3_add_63_U1_14 ( .A(fracta[14]), .B(fractb[14]), .CI(
        u3_add_63_carry[14]), .CO(u3_add_63_carry[15]), .S(u3_N17) );
  FA_X1 u3_add_63_U1_15 ( .A(fracta[15]), .B(fractb[15]), .CI(
        u3_add_63_carry[15]), .CO(u3_add_63_carry[16]), .S(u3_N18) );
  FA_X1 u3_add_63_U1_16 ( .A(fracta[16]), .B(fractb[16]), .CI(
        u3_add_63_carry[16]), .CO(u3_add_63_carry[17]), .S(u3_N19) );
  FA_X1 u3_add_63_U1_17 ( .A(fracta[17]), .B(fractb[17]), .CI(
        u3_add_63_carry[17]), .CO(u3_add_63_carry[18]), .S(u3_N20) );
  FA_X1 u3_add_63_U1_18 ( .A(fracta[18]), .B(fractb[18]), .CI(
        u3_add_63_carry[18]), .CO(u3_add_63_carry[19]), .S(u3_N21) );
  FA_X1 u3_add_63_U1_19 ( .A(fracta[19]), .B(fractb[19]), .CI(
        u3_add_63_carry[19]), .CO(u3_add_63_carry[20]), .S(u3_N22) );
  FA_X1 u3_add_63_U1_20 ( .A(fracta[20]), .B(fractb[20]), .CI(
        u3_add_63_carry[20]), .CO(u3_add_63_carry[21]), .S(u3_N23) );
  FA_X1 u3_add_63_U1_21 ( .A(fracta[21]), .B(fractb[21]), .CI(
        u3_add_63_carry[21]), .CO(u3_add_63_carry[22]), .S(u3_N24) );
  FA_X1 u3_add_63_U1_22 ( .A(fracta[22]), .B(fractb[22]), .CI(
        u3_add_63_carry[22]), .CO(u3_add_63_carry[23]), .S(u3_N25) );
  FA_X1 u3_add_63_U1_23 ( .A(fracta[23]), .B(fractb[23]), .CI(
        u3_add_63_carry[23]), .CO(u3_add_63_carry[24]), .S(u3_N26) );
  FA_X1 u3_add_63_U1_24 ( .A(fracta[24]), .B(fractb[24]), .CI(
        u3_add_63_carry[24]), .CO(u3_add_63_carry[25]), .S(u3_N27) );
  FA_X1 u3_add_63_U1_25 ( .A(fracta[25]), .B(fractb[25]), .CI(
        u3_add_63_carry[25]), .CO(u3_add_63_carry[26]), .S(u3_N28) );
  FA_X1 u3_add_63_U1_26 ( .A(fracta[26]), .B(fractb[26]), .CI(
        u3_add_63_carry[26]), .CO(u3_add_63_carry[27]), .S(u3_N29) );
  FA_X1 u3_add_63_U1_27 ( .A(fracta[27]), .B(fractb[27]), .CI(
        u3_add_63_carry[27]), .CO(u3_add_63_carry[28]), .S(u3_N30) );
  FA_X1 u3_add_63_U1_28 ( .A(fracta[28]), .B(fractb[28]), .CI(
        u3_add_63_carry[28]), .CO(u3_add_63_carry[29]), .S(u3_N31) );
  FA_X1 u3_add_63_U1_29 ( .A(fracta[29]), .B(fractb[29]), .CI(
        u3_add_63_carry[29]), .CO(u3_add_63_carry[30]), .S(u3_N32) );
  FA_X1 u3_add_63_U1_30 ( .A(fracta[30]), .B(fractb[30]), .CI(
        u3_add_63_carry[30]), .CO(u3_add_63_carry[31]), .S(u3_N33) );
  FA_X1 u3_add_63_U1_31 ( .A(fracta[31]), .B(fractb[31]), .CI(
        u3_add_63_carry[31]), .CO(u3_add_63_carry[32]), .S(u3_N34) );
  FA_X1 u3_add_63_U1_32 ( .A(fracta[32]), .B(fractb[32]), .CI(
        u3_add_63_carry[32]), .CO(u3_add_63_carry[33]), .S(u3_N35) );
  FA_X1 u3_add_63_U1_33 ( .A(fracta[33]), .B(fractb[33]), .CI(
        u3_add_63_carry[33]), .CO(u3_add_63_carry[34]), .S(u3_N36) );
  FA_X1 u3_add_63_U1_34 ( .A(fracta[34]), .B(fractb[34]), .CI(
        u3_add_63_carry[34]), .CO(u3_add_63_carry[35]), .S(u3_N37) );
  FA_X1 u3_add_63_U1_35 ( .A(fracta[35]), .B(fractb[35]), .CI(
        u3_add_63_carry[35]), .CO(u3_add_63_carry[36]), .S(u3_N38) );
  FA_X1 u3_add_63_U1_36 ( .A(fracta[36]), .B(fractb[36]), .CI(
        u3_add_63_carry[36]), .CO(u3_add_63_carry[37]), .S(u3_N39) );
  FA_X1 u3_add_63_U1_37 ( .A(fracta[37]), .B(fractb[37]), .CI(
        u3_add_63_carry[37]), .CO(u3_add_63_carry[38]), .S(u3_N40) );
  FA_X1 u3_add_63_U1_38 ( .A(fracta[38]), .B(fractb[38]), .CI(
        u3_add_63_carry[38]), .CO(u3_add_63_carry[39]), .S(u3_N41) );
  FA_X1 u3_add_63_U1_39 ( .A(fracta[39]), .B(fractb[39]), .CI(
        u3_add_63_carry[39]), .CO(u3_add_63_carry[40]), .S(u3_N42) );
  FA_X1 u3_add_63_U1_40 ( .A(fracta[40]), .B(fractb[40]), .CI(
        u3_add_63_carry[40]), .CO(u3_add_63_carry[41]), .S(u3_N43) );
  FA_X1 u3_add_63_U1_41 ( .A(fracta[41]), .B(fractb[41]), .CI(
        u3_add_63_carry[41]), .CO(u3_add_63_carry[42]), .S(u3_N44) );
  FA_X1 u3_add_63_U1_42 ( .A(fracta[42]), .B(fractb[42]), .CI(
        u3_add_63_carry[42]), .CO(u3_add_63_carry[43]), .S(u3_N45) );
  FA_X1 u3_add_63_U1_43 ( .A(fracta[43]), .B(fractb[43]), .CI(
        u3_add_63_carry[43]), .CO(u3_add_63_carry[44]), .S(u3_N46) );
  FA_X1 u3_add_63_U1_44 ( .A(fracta[44]), .B(fractb[44]), .CI(
        u3_add_63_carry[44]), .CO(u3_add_63_carry[45]), .S(u3_N47) );
  FA_X1 u3_add_63_U1_45 ( .A(fracta[45]), .B(fractb[45]), .CI(
        u3_add_63_carry[45]), .CO(u3_add_63_carry[46]), .S(u3_N48) );
  FA_X1 u3_add_63_U1_46 ( .A(fracta[46]), .B(fractb[46]), .CI(
        u3_add_63_carry[46]), .CO(u3_add_63_carry[47]), .S(u3_N49) );
  FA_X1 u3_add_63_U1_47 ( .A(fracta[47]), .B(fractb[47]), .CI(
        u3_add_63_carry[47]), .CO(u3_add_63_carry[48]), .S(u3_N50) );
  FA_X1 u3_add_63_U1_48 ( .A(fracta[48]), .B(fractb[48]), .CI(
        u3_add_63_carry[48]), .CO(u3_add_63_carry[49]), .S(u3_N51) );
  FA_X1 u3_add_63_U1_49 ( .A(fracta[49]), .B(fractb[49]), .CI(
        u3_add_63_carry[49]), .CO(u3_add_63_carry[50]), .S(u3_N52) );
  FA_X1 u3_add_63_U1_50 ( .A(fracta[50]), .B(fractb[50]), .CI(
        u3_add_63_carry[50]), .CO(u3_add_63_carry[51]), .S(u3_N53) );
  FA_X1 u3_add_63_U1_51 ( .A(fracta[51]), .B(fractb[51]), .CI(
        u3_add_63_carry[51]), .CO(u3_add_63_carry[52]), .S(u3_N54) );
  FA_X1 u3_add_63_U1_52 ( .A(fracta[52]), .B(fractb[52]), .CI(
        u3_add_63_carry[52]), .CO(u3_add_63_carry[53]), .S(u3_N55) );
  FA_X1 u3_add_63_U1_53 ( .A(fracta[53]), .B(fractb[53]), .CI(
        u3_add_63_carry[53]), .CO(u3_add_63_carry[54]), .S(u3_N56) );
  FA_X1 u3_add_63_U1_54 ( .A(fracta[54]), .B(fractb[54]), .CI(
        u3_add_63_carry[54]), .CO(u3_add_63_carry[55]), .S(u3_N57) );
  FA_X1 u3_add_63_U1_55 ( .A(fracta[55]), .B(fractb[55]), .CI(
        u3_add_63_carry[55]), .CO(u3_N59), .S(u3_N58) );
  XOR2_X1 u2_add_120_U2 ( .A(u2_add_120_carry[10]), .B(u2_exp_tmp4_10_), .Z(
        u2_N64) );
  INV_X4 u2_add_120_U1 ( .A(n2800), .ZN(u2_N54) );
  HA_X1 u2_add_120_U1_1_1 ( .A(u2_exp_tmp4_1_), .B(n2800), .CO(
        u2_add_120_carry[2]), .S(u2_N55) );
  HA_X1 u2_add_120_U1_1_2 ( .A(u2_exp_tmp4_2_), .B(u2_add_120_carry[2]), .CO(
        u2_add_120_carry[3]), .S(u2_N56) );
  HA_X1 u2_add_120_U1_1_3 ( .A(u2_exp_tmp4_3_), .B(u2_add_120_carry[3]), .CO(
        u2_add_120_carry[4]), .S(u2_N57) );
  HA_X1 u2_add_120_U1_1_4 ( .A(u2_exp_tmp4_4_), .B(u2_add_120_carry[4]), .CO(
        u2_add_120_carry[5]), .S(u2_N58) );
  HA_X1 u2_add_120_U1_1_5 ( .A(n2799), .B(u2_add_120_carry[5]), .CO(
        u2_add_120_carry[6]), .S(u2_N59) );
  HA_X1 u2_add_120_U1_1_6 ( .A(n2798), .B(u2_add_120_carry[6]), .CO(
        u2_add_120_carry[7]), .S(u2_N60) );
  HA_X1 u2_add_120_U1_1_7 ( .A(n2797), .B(u2_add_120_carry[7]), .CO(
        u2_add_120_carry[8]), .S(u2_N61) );
  HA_X1 u2_add_120_U1_1_8 ( .A(n2796), .B(u2_add_120_carry[8]), .CO(
        u2_add_120_carry[9]), .S(u2_N62) );
  HA_X1 u2_add_120_U1_1_9 ( .A(n2795), .B(u2_add_120_carry[9]), .CO(
        u2_add_120_carry[10]), .S(u2_N63) );
  XOR2_X1 u2_add_118_U2 ( .A(u2_add_118_carry[10]), .B(n6016), .Z(
        u2_exp_tmp3_10_) );
  INV_X4 u2_add_118_U1 ( .A(n6031), .ZN(u2_exp_tmp3_0_) );
  HA_X1 u2_add_118_U1_1_1 ( .A(n6029), .B(n6031), .CO(u2_add_118_carry[2]), 
        .S(u2_exp_tmp3_1_) );
  HA_X1 u2_add_118_U1_1_2 ( .A(n6027), .B(u2_add_118_carry[2]), .CO(
        u2_add_118_carry[3]), .S(u2_exp_tmp3_2_) );
  HA_X1 u2_add_118_U1_1_3 ( .A(n6025), .B(u2_add_118_carry[3]), .CO(
        u2_add_118_carry[4]), .S(u2_exp_tmp3_3_) );
  HA_X1 u2_add_118_U1_1_4 ( .A(n6023), .B(u2_add_118_carry[4]), .CO(
        u2_add_118_carry[5]), .S(u2_exp_tmp3_4_) );
  HA_X1 u2_add_118_U1_1_5 ( .A(n6022), .B(u2_add_118_carry[5]), .CO(
        u2_add_118_carry[6]), .S(u2_exp_tmp3_5_) );
  HA_X1 u2_add_118_U1_1_6 ( .A(n6021), .B(u2_add_118_carry[6]), .CO(
        u2_add_118_carry[7]), .S(u2_exp_tmp3_6_) );
  HA_X1 u2_add_118_U1_1_7 ( .A(n6020), .B(u2_add_118_carry[7]), .CO(
        u2_add_118_carry[8]), .S(u2_exp_tmp3_7_) );
  HA_X1 u2_add_118_U1_1_8 ( .A(n6019), .B(u2_add_118_carry[8]), .CO(
        u2_add_118_carry[9]), .S(u2_exp_tmp3_8_) );
  HA_X1 u2_add_118_U1_1_9 ( .A(n6018), .B(u2_add_118_carry[9]), .CO(
        u2_add_118_carry[10]), .S(u2_exp_tmp3_9_) );
  AND2_X4 u2_add_115_U2 ( .A1(opb_r[52]), .A2(opa_r[52]), .ZN(u2_add_115_n2)
         );
  XOR2_X2 u2_add_115_U1 ( .A(opb_r[52]), .B(opa_r[52]), .Z(u2_N18) );
  FA_X1 u2_add_115_U1_1 ( .A(opa_r[53]), .B(opb_r[53]), .CI(u2_add_115_n2), 
        .CO(u2_add_115_carry[2]), .S(u2_N19) );
  FA_X1 u2_add_115_U1_2 ( .A(opa_r[54]), .B(opb_r[54]), .CI(
        u2_add_115_carry[2]), .CO(u2_add_115_carry[3]), .S(u2_N20) );
  FA_X1 u2_add_115_U1_3 ( .A(opa_r[55]), .B(opb_r[55]), .CI(
        u2_add_115_carry[3]), .CO(u2_add_115_carry[4]), .S(u2_N21) );
  FA_X1 u2_add_115_U1_4 ( .A(opa_r[56]), .B(opb_r[56]), .CI(
        u2_add_115_carry[4]), .CO(u2_add_115_carry[5]), .S(u2_N22) );
  FA_X1 u2_add_115_U1_5 ( .A(opa_r[57]), .B(opb_r[57]), .CI(
        u2_add_115_carry[5]), .CO(u2_add_115_carry[6]), .S(u2_N23) );
  FA_X1 u2_add_115_U1_6 ( .A(opa_r[58]), .B(opb_r[58]), .CI(
        u2_add_115_carry[6]), .CO(u2_add_115_carry[7]), .S(u2_N24) );
  FA_X1 u2_add_115_U1_7 ( .A(opa_r[59]), .B(opb_r[59]), .CI(
        u2_add_115_carry[7]), .CO(u2_add_115_carry[8]), .S(u2_N25) );
  FA_X1 u2_add_115_U1_8 ( .A(opa_r[60]), .B(opb_r[60]), .CI(
        u2_add_115_carry[8]), .CO(u2_add_115_carry[9]), .S(u2_N26) );
  FA_X1 u2_add_115_U1_9 ( .A(opa_r[61]), .B(opb_r[61]), .CI(
        u2_add_115_carry[9]), .CO(u2_add_115_carry[10]), .S(u2_N27) );
  FA_X1 u2_add_115_U1_10 ( .A(opa_r[62]), .B(opb_r[62]), .CI(
        u2_add_115_carry[10]), .CO(u2_N29), .S(u2_N28) );
  INV_X4 u2_sub_115_U15 ( .A(opb_r[52]), .ZN(u2_sub_115_n13) );
  INV_X4 u2_sub_115_U14 ( .A(opb_r[53]), .ZN(u2_sub_115_n12) );
  INV_X4 u2_sub_115_U13 ( .A(opb_r[54]), .ZN(u2_sub_115_n11) );
  INV_X4 u2_sub_115_U12 ( .A(opb_r[55]), .ZN(u2_sub_115_n10) );
  INV_X4 u2_sub_115_U11 ( .A(opb_r[56]), .ZN(u2_sub_115_n9) );
  INV_X4 u2_sub_115_U10 ( .A(opb_r[57]), .ZN(u2_sub_115_n8) );
  INV_X4 u2_sub_115_U9 ( .A(opb_r[58]), .ZN(u2_sub_115_n7) );
  INV_X4 u2_sub_115_U8 ( .A(opb_r[59]), .ZN(u2_sub_115_n6) );
  INV_X4 u2_sub_115_U7 ( .A(opb_r[60]), .ZN(u2_sub_115_n5) );
  INV_X4 u2_sub_115_U6 ( .A(opb_r[61]), .ZN(u2_sub_115_n4) );
  INV_X4 u2_sub_115_U5 ( .A(opb_r[62]), .ZN(u2_sub_115_n3) );
  INV_X4 u2_sub_115_U4 ( .A(u2_sub_115_carry[11]), .ZN(u2_N17) );
  INV_X4 u2_sub_115_U3 ( .A(opa_r[52]), .ZN(u2_sub_115_n1) );
  XNOR2_X2 u2_sub_115_U2 ( .A(u2_sub_115_n13), .B(opa_r[52]), .ZN(u2_N6) );
  NAND2_X2 u2_sub_115_U1 ( .A1(opb_r[52]), .A2(u2_sub_115_n1), .ZN(
        u2_sub_115_carry[1]) );
  FA_X1 u2_sub_115_U2_1 ( .A(opa_r[53]), .B(u2_sub_115_n12), .CI(
        u2_sub_115_carry[1]), .CO(u2_sub_115_carry[2]), .S(u2_N7) );
  FA_X1 u2_sub_115_U2_2 ( .A(opa_r[54]), .B(u2_sub_115_n11), .CI(
        u2_sub_115_carry[2]), .CO(u2_sub_115_carry[3]), .S(u2_N8) );
  FA_X1 u2_sub_115_U2_3 ( .A(opa_r[55]), .B(u2_sub_115_n10), .CI(
        u2_sub_115_carry[3]), .CO(u2_sub_115_carry[4]), .S(u2_N9) );
  FA_X1 u2_sub_115_U2_4 ( .A(opa_r[56]), .B(u2_sub_115_n9), .CI(
        u2_sub_115_carry[4]), .CO(u2_sub_115_carry[5]), .S(u2_N10) );
  FA_X1 u2_sub_115_U2_5 ( .A(opa_r[57]), .B(u2_sub_115_n8), .CI(
        u2_sub_115_carry[5]), .CO(u2_sub_115_carry[6]), .S(u2_N11) );
  FA_X1 u2_sub_115_U2_6 ( .A(opa_r[58]), .B(u2_sub_115_n7), .CI(
        u2_sub_115_carry[6]), .CO(u2_sub_115_carry[7]), .S(u2_N12) );
  FA_X1 u2_sub_115_U2_7 ( .A(opa_r[59]), .B(u2_sub_115_n6), .CI(
        u2_sub_115_carry[7]), .CO(u2_sub_115_carry[8]), .S(u2_N13) );
  FA_X1 u2_sub_115_U2_8 ( .A(opa_r[60]), .B(u2_sub_115_n5), .CI(
        u2_sub_115_carry[8]), .CO(u2_sub_115_carry[9]), .S(u2_N14) );
  FA_X1 u2_sub_115_U2_9 ( .A(opa_r[61]), .B(u2_sub_115_n4), .CI(
        u2_sub_115_carry[9]), .CO(u2_sub_115_carry[10]), .S(u2_N15) );
  FA_X1 u2_sub_115_U2_10 ( .A(opa_r[62]), .B(u2_sub_115_n3), .CI(
        u2_sub_115_carry[10]), .CO(u2_sub_115_carry[11]), .S(u2_N16) );
  NOR2_X1 u1_gt_239_U168 ( .A1(n6159), .A2(u1_gt_239_n7), .ZN(u1_gt_239_n112)
         );
  NOR2_X1 u1_gt_239_U167 ( .A1(u1_gt_239_n109), .A2(n6208), .ZN(u1_gt_239_n167) );
  AOI21_X1 u1_gt_239_U166 ( .B1(u1_gt_239_n167), .B2(u1_gt_239_n97), .A(n6210), 
        .ZN(u1_gt_239_n166) );
  AOI221_X1 u1_gt_239_U165 ( .B1(n6186), .B2(u1_gt_239_n110), .C1(n6197), .C2(
        u1_gt_239_n108), .A(u1_gt_239_n166), .ZN(u1_gt_239_n165) );
  AOI221_X1 u1_gt_239_U164 ( .B1(n6122), .B2(u1_gt_239_n75), .C1(n6211), .C2(
        u1_gt_239_n86), .A(u1_gt_239_n165), .ZN(u1_gt_239_n164) );
  AOI221_X1 u1_gt_239_U163 ( .B1(n6164), .B2(u1_gt_239_n12), .C1(n6175), .C2(
        u1_gt_239_n23), .A(u1_gt_239_n164), .ZN(u1_gt_239_n163) );
  AOI221_X1 u1_gt_239_U162 ( .B1(n6104), .B2(u1_gt_239_n58), .C1(n6111), .C2(
        u1_gt_239_n64), .A(u1_gt_239_n163), .ZN(u1_gt_239_n162) );
  AOI221_X1 u1_gt_239_U161 ( .B1(n6156), .B2(u1_gt_239_n4), .C1(n6157), .C2(
        u1_gt_239_n5), .A(u1_gt_239_n162), .ZN(u1_gt_239_n161) );
  AOI221_X1 u1_gt_239_U160 ( .B1(n6102), .B2(u1_gt_239_n56), .C1(n6103), .C2(
        u1_gt_239_n57), .A(u1_gt_239_n161), .ZN(u1_gt_239_n160) );
  AOI221_X1 u1_gt_239_U159 ( .B1(n6154), .B2(u1_gt_239_n2), .C1(n6155), .C2(
        u1_gt_239_n3), .A(u1_gt_239_n160), .ZN(u1_gt_239_n159) );
  AOI221_X1 u1_gt_239_U158 ( .B1(n6100), .B2(u1_gt_239_n54), .C1(n6101), .C2(
        u1_gt_239_n55), .A(u1_gt_239_n159), .ZN(u1_gt_239_n158) );
  AOI221_X1 u1_gt_239_U157 ( .B1(n6153), .B2(u1_gt_239_n1), .C1(n6207), .C2(
        u1_gt_239_n53), .A(u1_gt_239_n158), .ZN(u1_gt_239_n157) );
  AOI221_X1 u1_gt_239_U156 ( .B1(n6151), .B2(u1_gt_239_n106), .C1(n6152), .C2(
        u1_gt_239_n107), .A(u1_gt_239_n157), .ZN(u1_gt_239_n156) );
  AOI221_X1 u1_gt_239_U155 ( .B1(n6205), .B2(u1_gt_239_n51), .C1(n6206), .C2(
        u1_gt_239_n52), .A(u1_gt_239_n156), .ZN(u1_gt_239_n155) );
  AOI221_X1 u1_gt_239_U154 ( .B1(n6149), .B2(u1_gt_239_n104), .C1(n6150), .C2(
        u1_gt_239_n105), .A(u1_gt_239_n155), .ZN(u1_gt_239_n154) );
  AOI221_X1 u1_gt_239_U153 ( .B1(n6203), .B2(u1_gt_239_n49), .C1(n6204), .C2(
        u1_gt_239_n50), .A(u1_gt_239_n154), .ZN(u1_gt_239_n153) );
  AOI221_X1 u1_gt_239_U152 ( .B1(n6147), .B2(u1_gt_239_n102), .C1(n6148), .C2(
        u1_gt_239_n103), .A(u1_gt_239_n153), .ZN(u1_gt_239_n152) );
  AOI221_X1 u1_gt_239_U151 ( .B1(n6201), .B2(u1_gt_239_n47), .C1(n6202), .C2(
        u1_gt_239_n48), .A(u1_gt_239_n152), .ZN(u1_gt_239_n151) );
  AOI221_X1 u1_gt_239_U150 ( .B1(n6145), .B2(u1_gt_239_n100), .C1(n6146), .C2(
        u1_gt_239_n101), .A(u1_gt_239_n151), .ZN(u1_gt_239_n150) );
  AOI221_X1 u1_gt_239_U149 ( .B1(n6199), .B2(u1_gt_239_n45), .C1(n6200), .C2(
        u1_gt_239_n46), .A(u1_gt_239_n150), .ZN(u1_gt_239_n149) );
  AOI221_X1 u1_gt_239_U148 ( .B1(n6143), .B2(u1_gt_239_n98), .C1(n6144), .C2(
        u1_gt_239_n99), .A(u1_gt_239_n149), .ZN(u1_gt_239_n148) );
  AOI221_X1 u1_gt_239_U147 ( .B1(n6196), .B2(u1_gt_239_n43), .C1(n6198), .C2(
        u1_gt_239_n44), .A(u1_gt_239_n148), .ZN(u1_gt_239_n147) );
  AOI221_X1 u1_gt_239_U146 ( .B1(n6141), .B2(u1_gt_239_n95), .C1(n6142), .C2(
        u1_gt_239_n96), .A(u1_gt_239_n147), .ZN(u1_gt_239_n146) );
  AOI221_X1 u1_gt_239_U145 ( .B1(n6194), .B2(u1_gt_239_n41), .C1(n6195), .C2(
        u1_gt_239_n42), .A(u1_gt_239_n146), .ZN(u1_gt_239_n145) );
  AOI221_X1 u1_gt_239_U144 ( .B1(n6139), .B2(u1_gt_239_n93), .C1(n6140), .C2(
        u1_gt_239_n94), .A(u1_gt_239_n145), .ZN(u1_gt_239_n144) );
  AOI221_X1 u1_gt_239_U143 ( .B1(n6192), .B2(u1_gt_239_n39), .C1(n6193), .C2(
        u1_gt_239_n40), .A(u1_gt_239_n144), .ZN(u1_gt_239_n143) );
  AOI221_X1 u1_gt_239_U142 ( .B1(n6137), .B2(u1_gt_239_n91), .C1(n6138), .C2(
        u1_gt_239_n92), .A(u1_gt_239_n143), .ZN(u1_gt_239_n142) );
  AOI221_X1 u1_gt_239_U141 ( .B1(n6190), .B2(u1_gt_239_n37), .C1(n6191), .C2(
        u1_gt_239_n38), .A(u1_gt_239_n142), .ZN(u1_gt_239_n141) );
  AOI221_X1 u1_gt_239_U140 ( .B1(n6135), .B2(u1_gt_239_n89), .C1(n6136), .C2(
        u1_gt_239_n90), .A(u1_gt_239_n141), .ZN(u1_gt_239_n140) );
  AOI221_X1 u1_gt_239_U139 ( .B1(n6188), .B2(u1_gt_239_n35), .C1(n6189), .C2(
        u1_gt_239_n36), .A(u1_gt_239_n140), .ZN(u1_gt_239_n139) );
  AOI221_X1 u1_gt_239_U138 ( .B1(n6133), .B2(u1_gt_239_n87), .C1(n6134), .C2(
        u1_gt_239_n88), .A(u1_gt_239_n139), .ZN(u1_gt_239_n138) );
  AOI221_X1 u1_gt_239_U137 ( .B1(n6185), .B2(u1_gt_239_n33), .C1(n6187), .C2(
        u1_gt_239_n34), .A(u1_gt_239_n138), .ZN(u1_gt_239_n137) );
  AOI221_X1 u1_gt_239_U136 ( .B1(n6131), .B2(u1_gt_239_n84), .C1(n6132), .C2(
        u1_gt_239_n85), .A(u1_gt_239_n137), .ZN(u1_gt_239_n136) );
  AOI221_X1 u1_gt_239_U135 ( .B1(n6183), .B2(u1_gt_239_n31), .C1(n6184), .C2(
        u1_gt_239_n32), .A(u1_gt_239_n136), .ZN(u1_gt_239_n135) );
  AOI221_X1 u1_gt_239_U134 ( .B1(n6129), .B2(u1_gt_239_n82), .C1(n6130), .C2(
        u1_gt_239_n83), .A(u1_gt_239_n135), .ZN(u1_gt_239_n134) );
  AOI221_X1 u1_gt_239_U133 ( .B1(n6181), .B2(u1_gt_239_n29), .C1(n6182), .C2(
        u1_gt_239_n30), .A(u1_gt_239_n134), .ZN(u1_gt_239_n133) );
  AOI221_X1 u1_gt_239_U132 ( .B1(n6127), .B2(u1_gt_239_n80), .C1(n6128), .C2(
        u1_gt_239_n81), .A(u1_gt_239_n133), .ZN(u1_gt_239_n132) );
  AOI221_X1 u1_gt_239_U131 ( .B1(n6179), .B2(u1_gt_239_n27), .C1(n6180), .C2(
        u1_gt_239_n28), .A(u1_gt_239_n132), .ZN(u1_gt_239_n131) );
  AOI221_X1 u1_gt_239_U130 ( .B1(n6125), .B2(u1_gt_239_n78), .C1(n6126), .C2(
        u1_gt_239_n79), .A(u1_gt_239_n131), .ZN(u1_gt_239_n130) );
  AOI221_X1 u1_gt_239_U129 ( .B1(n6177), .B2(u1_gt_239_n25), .C1(n6178), .C2(
        u1_gt_239_n26), .A(u1_gt_239_n130), .ZN(u1_gt_239_n129) );
  AOI221_X1 u1_gt_239_U128 ( .B1(n6123), .B2(u1_gt_239_n76), .C1(n6124), .C2(
        u1_gt_239_n77), .A(u1_gt_239_n129), .ZN(u1_gt_239_n128) );
  AOI221_X1 u1_gt_239_U127 ( .B1(n6174), .B2(u1_gt_239_n22), .C1(n6176), .C2(
        u1_gt_239_n24), .A(u1_gt_239_n128), .ZN(u1_gt_239_n127) );
  AOI221_X1 u1_gt_239_U126 ( .B1(n6120), .B2(u1_gt_239_n73), .C1(n6121), .C2(
        u1_gt_239_n74), .A(u1_gt_239_n127), .ZN(u1_gt_239_n126) );
  AOI221_X1 u1_gt_239_U125 ( .B1(n6172), .B2(u1_gt_239_n20), .C1(n6173), .C2(
        u1_gt_239_n21), .A(u1_gt_239_n126), .ZN(u1_gt_239_n125) );
  AOI221_X1 u1_gt_239_U124 ( .B1(n6118), .B2(u1_gt_239_n71), .C1(n6119), .C2(
        u1_gt_239_n72), .A(u1_gt_239_n125), .ZN(u1_gt_239_n124) );
  AOI221_X1 u1_gt_239_U123 ( .B1(n6170), .B2(u1_gt_239_n18), .C1(n6171), .C2(
        u1_gt_239_n19), .A(u1_gt_239_n124), .ZN(u1_gt_239_n123) );
  AOI221_X1 u1_gt_239_U122 ( .B1(n6116), .B2(u1_gt_239_n69), .C1(n6117), .C2(
        u1_gt_239_n70), .A(u1_gt_239_n123), .ZN(u1_gt_239_n122) );
  AOI221_X1 u1_gt_239_U121 ( .B1(n6168), .B2(u1_gt_239_n16), .C1(n6169), .C2(
        u1_gt_239_n17), .A(u1_gt_239_n122), .ZN(u1_gt_239_n121) );
  AOI221_X1 u1_gt_239_U120 ( .B1(n6114), .B2(u1_gt_239_n67), .C1(n6115), .C2(
        u1_gt_239_n68), .A(u1_gt_239_n121), .ZN(u1_gt_239_n120) );
  AOI221_X1 u1_gt_239_U119 ( .B1(n6166), .B2(u1_gt_239_n14), .C1(n6167), .C2(
        u1_gt_239_n15), .A(u1_gt_239_n120), .ZN(u1_gt_239_n119) );
  AOI221_X1 u1_gt_239_U118 ( .B1(n6112), .B2(u1_gt_239_n65), .C1(n6113), .C2(
        u1_gt_239_n66), .A(u1_gt_239_n119), .ZN(u1_gt_239_n118) );
  AOI221_X1 u1_gt_239_U117 ( .B1(n6163), .B2(u1_gt_239_n11), .C1(n6165), .C2(
        u1_gt_239_n13), .A(u1_gt_239_n118), .ZN(u1_gt_239_n117) );
  AOI221_X1 u1_gt_239_U116 ( .B1(n6109), .B2(u1_gt_239_n62), .C1(n6110), .C2(
        u1_gt_239_n63), .A(u1_gt_239_n117), .ZN(u1_gt_239_n116) );
  AOI221_X1 u1_gt_239_U115 ( .B1(n6161), .B2(u1_gt_239_n9), .C1(n6162), .C2(
        u1_gt_239_n10), .A(u1_gt_239_n116), .ZN(u1_gt_239_n115) );
  AOI221_X1 u1_gt_239_U114 ( .B1(n6107), .B2(u1_gt_239_n60), .C1(n6108), .C2(
        u1_gt_239_n61), .A(u1_gt_239_n115), .ZN(u1_gt_239_n114) );
  AOI221_X1 u1_gt_239_U113 ( .B1(n6159), .B2(u1_gt_239_n7), .C1(n6160), .C2(
        u1_gt_239_n8), .A(u1_gt_239_n114), .ZN(u1_gt_239_n113) );
  OAI22_X1 u1_gt_239_U112 ( .A1(u1_gt_239_n112), .A2(u1_gt_239_n113), .B1(
        n6105), .B2(u1_gt_239_n59), .ZN(u1_gt_239_n111) );
  OAI21_X1 u1_gt_239_U111 ( .B1(n6158), .B2(u1_gt_239_n6), .A(u1_gt_239_n111), 
        .ZN(u1_fractb_lt_fracta) );
  INV_X4 u1_gt_239_U110 ( .A(n6211), .ZN(u1_gt_239_n110) );
  INV_X4 u1_gt_239_U109 ( .A(n6209), .ZN(u1_gt_239_n109) );
  INV_X4 u1_gt_239_U108 ( .A(u1_gt_239_n167), .ZN(u1_gt_239_n108) );
  INV_X4 u1_gt_239_U107 ( .A(n6207), .ZN(u1_gt_239_n107) );
  INV_X4 u1_gt_239_U106 ( .A(n6206), .ZN(u1_gt_239_n106) );
  INV_X4 u1_gt_239_U105 ( .A(n6205), .ZN(u1_gt_239_n105) );
  INV_X4 u1_gt_239_U104 ( .A(n6204), .ZN(u1_gt_239_n104) );
  INV_X4 u1_gt_239_U103 ( .A(n6203), .ZN(u1_gt_239_n103) );
  INV_X4 u1_gt_239_U102 ( .A(n6202), .ZN(u1_gt_239_n102) );
  INV_X4 u1_gt_239_U101 ( .A(n6201), .ZN(u1_gt_239_n101) );
  INV_X4 u1_gt_239_U100 ( .A(n6200), .ZN(u1_gt_239_n100) );
  INV_X4 u1_gt_239_U99 ( .A(n6199), .ZN(u1_gt_239_n99) );
  INV_X4 u1_gt_239_U98 ( .A(n6198), .ZN(u1_gt_239_n98) );
  INV_X4 u1_gt_239_U97 ( .A(n6197), .ZN(u1_gt_239_n97) );
  INV_X4 u1_gt_239_U96 ( .A(n6196), .ZN(u1_gt_239_n96) );
  INV_X4 u1_gt_239_U95 ( .A(n6195), .ZN(u1_gt_239_n95) );
  INV_X4 u1_gt_239_U94 ( .A(n6194), .ZN(u1_gt_239_n94) );
  INV_X4 u1_gt_239_U93 ( .A(n6193), .ZN(u1_gt_239_n93) );
  INV_X4 u1_gt_239_U92 ( .A(n6192), .ZN(u1_gt_239_n92) );
  INV_X4 u1_gt_239_U91 ( .A(n6191), .ZN(u1_gt_239_n91) );
  INV_X4 u1_gt_239_U90 ( .A(n6190), .ZN(u1_gt_239_n90) );
  INV_X4 u1_gt_239_U89 ( .A(n6189), .ZN(u1_gt_239_n89) );
  INV_X4 u1_gt_239_U88 ( .A(n6188), .ZN(u1_gt_239_n88) );
  INV_X4 u1_gt_239_U87 ( .A(n6187), .ZN(u1_gt_239_n87) );
  INV_X4 u1_gt_239_U86 ( .A(n6186), .ZN(u1_gt_239_n86) );
  INV_X4 u1_gt_239_U85 ( .A(n6185), .ZN(u1_gt_239_n85) );
  INV_X4 u1_gt_239_U84 ( .A(n6184), .ZN(u1_gt_239_n84) );
  INV_X4 u1_gt_239_U83 ( .A(n6183), .ZN(u1_gt_239_n83) );
  INV_X4 u1_gt_239_U82 ( .A(n6182), .ZN(u1_gt_239_n82) );
  INV_X4 u1_gt_239_U81 ( .A(n6181), .ZN(u1_gt_239_n81) );
  INV_X4 u1_gt_239_U80 ( .A(n6180), .ZN(u1_gt_239_n80) );
  INV_X4 u1_gt_239_U79 ( .A(n6179), .ZN(u1_gt_239_n79) );
  INV_X4 u1_gt_239_U78 ( .A(n6178), .ZN(u1_gt_239_n78) );
  INV_X4 u1_gt_239_U77 ( .A(n6177), .ZN(u1_gt_239_n77) );
  INV_X4 u1_gt_239_U76 ( .A(n6176), .ZN(u1_gt_239_n76) );
  INV_X4 u1_gt_239_U75 ( .A(n6175), .ZN(u1_gt_239_n75) );
  INV_X4 u1_gt_239_U74 ( .A(n6174), .ZN(u1_gt_239_n74) );
  INV_X4 u1_gt_239_U73 ( .A(n6173), .ZN(u1_gt_239_n73) );
  INV_X4 u1_gt_239_U72 ( .A(n6172), .ZN(u1_gt_239_n72) );
  INV_X4 u1_gt_239_U71 ( .A(n6171), .ZN(u1_gt_239_n71) );
  INV_X4 u1_gt_239_U70 ( .A(n6170), .ZN(u1_gt_239_n70) );
  INV_X4 u1_gt_239_U69 ( .A(n6169), .ZN(u1_gt_239_n69) );
  INV_X4 u1_gt_239_U68 ( .A(n6168), .ZN(u1_gt_239_n68) );
  INV_X4 u1_gt_239_U67 ( .A(n6167), .ZN(u1_gt_239_n67) );
  INV_X4 u1_gt_239_U66 ( .A(n6166), .ZN(u1_gt_239_n66) );
  INV_X4 u1_gt_239_U65 ( .A(n6165), .ZN(u1_gt_239_n65) );
  INV_X4 u1_gt_239_U64 ( .A(n6164), .ZN(u1_gt_239_n64) );
  INV_X4 u1_gt_239_U63 ( .A(n6163), .ZN(u1_gt_239_n63) );
  INV_X4 u1_gt_239_U62 ( .A(n6162), .ZN(u1_gt_239_n62) );
  INV_X4 u1_gt_239_U61 ( .A(n6161), .ZN(u1_gt_239_n61) );
  INV_X4 u1_gt_239_U60 ( .A(n6160), .ZN(u1_gt_239_n60) );
  INV_X4 u1_gt_239_U59 ( .A(n6158), .ZN(u1_gt_239_n59) );
  INV_X4 u1_gt_239_U58 ( .A(n6157), .ZN(u1_gt_239_n58) );
  INV_X4 u1_gt_239_U57 ( .A(n6156), .ZN(u1_gt_239_n57) );
  INV_X4 u1_gt_239_U56 ( .A(n6155), .ZN(u1_gt_239_n56) );
  INV_X4 u1_gt_239_U55 ( .A(n6154), .ZN(u1_gt_239_n55) );
  INV_X4 u1_gt_239_U54 ( .A(n6153), .ZN(u1_gt_239_n54) );
  INV_X4 u1_gt_239_U53 ( .A(n6152), .ZN(u1_gt_239_n53) );
  INV_X4 u1_gt_239_U52 ( .A(n6151), .ZN(u1_gt_239_n52) );
  INV_X4 u1_gt_239_U51 ( .A(n6150), .ZN(u1_gt_239_n51) );
  INV_X4 u1_gt_239_U50 ( .A(n6149), .ZN(u1_gt_239_n50) );
  INV_X4 u1_gt_239_U49 ( .A(n6148), .ZN(u1_gt_239_n49) );
  INV_X4 u1_gt_239_U48 ( .A(n6147), .ZN(u1_gt_239_n48) );
  INV_X4 u1_gt_239_U47 ( .A(n6146), .ZN(u1_gt_239_n47) );
  INV_X4 u1_gt_239_U46 ( .A(n6145), .ZN(u1_gt_239_n46) );
  INV_X4 u1_gt_239_U45 ( .A(n6144), .ZN(u1_gt_239_n45) );
  INV_X4 u1_gt_239_U44 ( .A(n6143), .ZN(u1_gt_239_n44) );
  INV_X4 u1_gt_239_U43 ( .A(n6142), .ZN(u1_gt_239_n43) );
  INV_X4 u1_gt_239_U42 ( .A(n6141), .ZN(u1_gt_239_n42) );
  INV_X4 u1_gt_239_U41 ( .A(n6140), .ZN(u1_gt_239_n41) );
  INV_X4 u1_gt_239_U40 ( .A(n6139), .ZN(u1_gt_239_n40) );
  INV_X4 u1_gt_239_U39 ( .A(n6138), .ZN(u1_gt_239_n39) );
  INV_X4 u1_gt_239_U38 ( .A(n6137), .ZN(u1_gt_239_n38) );
  INV_X4 u1_gt_239_U37 ( .A(n6136), .ZN(u1_gt_239_n37) );
  INV_X4 u1_gt_239_U36 ( .A(n6135), .ZN(u1_gt_239_n36) );
  INV_X4 u1_gt_239_U35 ( .A(n6134), .ZN(u1_gt_239_n35) );
  INV_X4 u1_gt_239_U34 ( .A(n6133), .ZN(u1_gt_239_n34) );
  INV_X4 u1_gt_239_U33 ( .A(n6132), .ZN(u1_gt_239_n33) );
  INV_X4 u1_gt_239_U32 ( .A(n6131), .ZN(u1_gt_239_n32) );
  INV_X4 u1_gt_239_U31 ( .A(n6130), .ZN(u1_gt_239_n31) );
  INV_X4 u1_gt_239_U30 ( .A(n6129), .ZN(u1_gt_239_n30) );
  INV_X4 u1_gt_239_U29 ( .A(n6128), .ZN(u1_gt_239_n29) );
  INV_X4 u1_gt_239_U28 ( .A(n6127), .ZN(u1_gt_239_n28) );
  INV_X4 u1_gt_239_U27 ( .A(n6126), .ZN(u1_gt_239_n27) );
  INV_X4 u1_gt_239_U26 ( .A(n6125), .ZN(u1_gt_239_n26) );
  INV_X4 u1_gt_239_U25 ( .A(n6124), .ZN(u1_gt_239_n25) );
  INV_X4 u1_gt_239_U24 ( .A(n6123), .ZN(u1_gt_239_n24) );
  INV_X4 u1_gt_239_U23 ( .A(n6122), .ZN(u1_gt_239_n23) );
  INV_X4 u1_gt_239_U22 ( .A(n6121), .ZN(u1_gt_239_n22) );
  INV_X4 u1_gt_239_U21 ( .A(n6120), .ZN(u1_gt_239_n21) );
  INV_X4 u1_gt_239_U20 ( .A(n6119), .ZN(u1_gt_239_n20) );
  INV_X4 u1_gt_239_U19 ( .A(n6118), .ZN(u1_gt_239_n19) );
  INV_X4 u1_gt_239_U18 ( .A(n6117), .ZN(u1_gt_239_n18) );
  INV_X4 u1_gt_239_U17 ( .A(n6116), .ZN(u1_gt_239_n17) );
  INV_X4 u1_gt_239_U16 ( .A(n6115), .ZN(u1_gt_239_n16) );
  INV_X4 u1_gt_239_U15 ( .A(n6114), .ZN(u1_gt_239_n15) );
  INV_X4 u1_gt_239_U14 ( .A(n6113), .ZN(u1_gt_239_n14) );
  INV_X4 u1_gt_239_U13 ( .A(n6112), .ZN(u1_gt_239_n13) );
  INV_X4 u1_gt_239_U12 ( .A(n6111), .ZN(u1_gt_239_n12) );
  INV_X4 u1_gt_239_U11 ( .A(n6110), .ZN(u1_gt_239_n11) );
  INV_X4 u1_gt_239_U10 ( .A(n6109), .ZN(u1_gt_239_n10) );
  INV_X4 u1_gt_239_U9 ( .A(n6108), .ZN(u1_gt_239_n9) );
  INV_X4 u1_gt_239_U8 ( .A(n6107), .ZN(u1_gt_239_n8) );
  INV_X4 u1_gt_239_U7 ( .A(n6106), .ZN(u1_gt_239_n7) );
  INV_X4 u1_gt_239_U6 ( .A(n6105), .ZN(u1_gt_239_n6) );
  INV_X4 u1_gt_239_U5 ( .A(n6104), .ZN(u1_gt_239_n5) );
  INV_X4 u1_gt_239_U4 ( .A(n6103), .ZN(u1_gt_239_n4) );
  INV_X4 u1_gt_239_U3 ( .A(n6102), .ZN(u1_gt_239_n3) );
  INV_X4 u1_gt_239_U2 ( .A(n6101), .ZN(u1_gt_239_n2) );
  INV_X4 u1_gt_239_U1 ( .A(n6100), .ZN(u1_gt_239_n1) );
  NOR2_X1 u1_srl_151_U418 ( .A1(u1_srl_151_n97), .A2(n6226), .ZN(
        u1_srl_151_n163) );
  AND2_X1 u1_srl_151_U417 ( .A1(n6221), .A2(n6222), .ZN(u1_srl_151_n198) );
  NOR2_X1 u1_srl_151_U416 ( .A1(n6222), .A2(n6221), .ZN(u1_srl_151_n199) );
  AOI22_X1 u1_srl_151_U415 ( .A1(u1_adj_op_28_), .A2(u1_srl_151_n15), .B1(
        n6253), .B2(u1_srl_151_n16), .ZN(u1_srl_151_n360) );
  OAI221_X1 u1_srl_151_U414 ( .B1(u1_srl_151_n6), .B2(u1_srl_151_n118), .C1(
        u1_srl_151_n12), .C2(u1_srl_151_n117), .A(u1_srl_151_n360), .ZN(
        u1_srl_151_n242) );
  AOI22_X1 u1_srl_151_U413 ( .A1(n6254), .A2(u1_srl_151_n15), .B1(
        u1_srl_151_n16), .B2(u1_adj_op_21_), .ZN(u1_srl_151_n359) );
  OAI221_X1 u1_srl_151_U412 ( .B1(u1_srl_151_n6), .B2(u1_srl_151_n122), .C1(
        u1_srl_151_n3), .C2(u1_srl_151_n121), .A(u1_srl_151_n359), .ZN(
        u1_srl_151_n243) );
  AOI22_X1 u1_srl_151_U411 ( .A1(u1_srl_151_n15), .A2(u1_adj_op_20_), .B1(
        u1_adj_op_17_), .B2(u1_srl_151_n16), .ZN(u1_srl_151_n358) );
  OAI221_X1 u1_srl_151_U410 ( .B1(u1_srl_151_n7), .B2(u1_srl_151_n127), .C1(
        u1_srl_151_n126), .C2(u1_srl_151_n3), .A(u1_srl_151_n358), .ZN(
        u1_srl_151_n153) );
  AOI22_X1 u1_srl_151_U409 ( .A1(u1_adj_op_16_), .A2(u1_srl_151_n15), .B1(
        n6260), .B2(u1_srl_151_n16), .ZN(u1_srl_151_n357) );
  OAI221_X1 u1_srl_151_U408 ( .B1(u1_srl_151_n7), .B2(u1_srl_151_n131), .C1(
        u1_srl_151_n3), .C2(u1_srl_151_n130), .A(u1_srl_151_n357), .ZN(
        u1_srl_151_n154) );
  AOI22_X1 u1_srl_151_U407 ( .A1(u1_srl_151_n10), .A2(u1_srl_151_n153), .B1(
        u1_srl_151_n2), .B2(u1_srl_151_n154), .ZN(u1_srl_151_n356) );
  AOI221_X1 u1_srl_151_U406 ( .B1(u1_srl_151_n242), .B2(u1_srl_151_n237), .C1(
        u1_srl_151_n243), .C2(u1_srl_151_n196), .A(u1_srl_151_n21), .ZN(
        u1_srl_151_n289) );
  AOI22_X1 u1_srl_151_U405 ( .A1(n6235), .A2(u1_srl_151_n15), .B1(n6256), .B2(
        u1_srl_151_n16), .ZN(u1_srl_151_n355) );
  OAI221_X1 u1_srl_151_U404 ( .B1(u1_srl_151_n7), .B2(u1_srl_151_n114), .C1(
        u1_srl_151_n12), .C2(u1_srl_151_n105), .A(u1_srl_151_n355), .ZN(
        u1_srl_151_n184) );
  AOI22_X1 u1_srl_151_U403 ( .A1(u1_adj_op_36_), .A2(u1_srl_151_n15), .B1(
        n6247), .B2(u1_srl_151_n16), .ZN(u1_srl_151_n354) );
  OAI221_X1 u1_srl_151_U402 ( .B1(u1_srl_151_n7), .B2(u1_srl_151_n109), .C1(
        u1_srl_151_n12), .C2(u1_srl_151_n108), .A(u1_srl_151_n354), .ZN(
        u1_srl_151_n245) );
  AOI22_X1 u1_srl_151_U401 ( .A1(u1_adj_op_32_), .A2(u1_srl_151_n15), .B1(
        n6251), .B2(u1_srl_151_n16), .ZN(u1_srl_151_n353) );
  OAI221_X1 u1_srl_151_U400 ( .B1(u1_srl_151_n7), .B2(u1_srl_151_n113), .C1(
        u1_srl_151_n12), .C2(u1_srl_151_n112), .A(u1_srl_151_n353), .ZN(
        u1_srl_151_n246) );
  AOI22_X1 u1_srl_151_U399 ( .A1(u1_adj_op_44_), .A2(u1_srl_151_n198), .B1(
        n6242), .B2(u1_srl_151_n199), .ZN(u1_srl_151_n352) );
  AOI221_X1 u1_srl_151_U398 ( .B1(u1_srl_151_n224), .B2(u1_adj_op_42_), .C1(
        u1_srl_151_n13), .C2(n6241), .A(u1_srl_151_n61), .ZN(u1_srl_151_n270)
         );
  AOI22_X1 u1_srl_151_U397 ( .A1(n6243), .A2(u1_srl_151_n198), .B1(
        u1_adj_op_37_), .B2(u1_srl_151_n199), .ZN(u1_srl_151_n351) );
  AOI221_X1 u1_srl_151_U396 ( .B1(u1_srl_151_n224), .B2(u1_adj_op_38_), .C1(
        u1_srl_151_n13), .C2(n6244), .A(u1_srl_151_n63), .ZN(u1_srl_151_n312)
         );
  OAI22_X1 u1_srl_151_U395 ( .A1(u1_srl_151_n58), .A2(u1_srl_151_n270), .B1(
        u1_srl_151_n5), .B2(u1_srl_151_n312), .ZN(u1_srl_151_n350) );
  AOI221_X1 u1_srl_151_U394 ( .B1(u1_srl_151_n245), .B2(u1_srl_151_n11), .C1(
        u1_srl_151_n246), .C2(u1_srl_151_n18), .A(u1_srl_151_n350), .ZN(
        u1_srl_151_n215) );
  AOI222_X1 u1_srl_151_U393 ( .A1(u1_srl_151_n163), .A2(u1_srl_151_n20), .B1(
        u1_srl_151_n139), .B2(u1_srl_151_n184), .C1(u1_srl_151_n145), .C2(
        u1_srl_151_n22), .ZN(u1_srl_151_n342) );
  NAND2_X1 u1_srl_151_U392 ( .A1(n6225), .A2(n6226), .ZN(u1_srl_151_n223) );
  AOI22_X1 u1_srl_151_U391 ( .A1(n6237), .A2(u1_srl_151_n15), .B1(n6240), .B2(
        u1_srl_151_n16), .ZN(u1_srl_151_n349) );
  AOI221_X1 u1_srl_151_U390 ( .B1(u1_srl_151_n224), .B2(n6239), .C1(
        u1_srl_151_n13), .C2(n6238), .A(u1_srl_151_n65), .ZN(u1_srl_151_n241)
         );
  AOI22_X1 u1_srl_151_U389 ( .A1(n4266), .A2(u1_srl_151_n15), .B1(n6236), .B2(
        u1_srl_151_n16), .ZN(u1_srl_151_n348) );
  AOI221_X1 u1_srl_151_U388 ( .B1(u1_srl_151_n224), .B2(n6234), .C1(
        u1_srl_151_n13), .C2(u1_adj_op_51_), .A(u1_srl_151_n67), .ZN(
        u1_srl_151_n179) );
  AOI22_X1 u1_srl_151_U387 ( .A1(u1_srl_151_n64), .A2(u1_srl_151_n18), .B1(
        u1_srl_151_n66), .B2(u1_srl_151_n11), .ZN(u1_srl_151_n187) );
  AOI22_X1 u1_srl_151_U386 ( .A1(n6230), .A2(u1_srl_151_n198), .B1(n6233), 
        .B2(u1_srl_151_n16), .ZN(u1_srl_151_n347) );
  OAI221_X1 u1_srl_151_U385 ( .B1(u1_srl_151_n7), .B2(u1_srl_151_n102), .C1(
        u1_srl_151_n12), .C2(u1_srl_151_n101), .A(u1_srl_151_n347), .ZN(
        u1_srl_151_n155) );
  AOI22_X1 u1_srl_151_U384 ( .A1(n6261), .A2(u1_srl_151_n198), .B1(n6229), 
        .B2(u1_srl_151_n16), .ZN(u1_srl_151_n346) );
  OAI221_X1 u1_srl_151_U383 ( .B1(u1_srl_151_n7), .B2(u1_srl_151_n135), .C1(
        u1_srl_151_n12), .C2(u1_srl_151_n134), .A(u1_srl_151_n346), .ZN(
        u1_srl_151_n152) );
  AOI22_X1 u1_srl_151_U382 ( .A1(u1_srl_151_n155), .A2(u1_srl_151_n143), .B1(
        u1_srl_151_n152), .B2(u1_srl_151_n141), .ZN(u1_srl_151_n344) );
  NAND3_X1 u1_srl_151_U381 ( .A1(u1_adj_op_0_), .A2(u1_srl_151_n15), .A3(
        u1_srl_151_n146), .ZN(u1_srl_151_n345) );
  OAI211_X1 u1_srl_151_U380 ( .C1(u1_srl_151_n223), .C2(u1_srl_151_n187), .A(
        u1_srl_151_n344), .B(u1_srl_151_n345), .ZN(u1_srl_151_n343) );
  NAND2_X1 u1_srl_151_U379 ( .A1(u1_srl_151_n342), .A2(u1_srl_151_n23), .ZN(
        u1_adj_op_out_sft_0_) );
  AOI22_X1 u1_srl_151_U378 ( .A1(n6249), .A2(u1_srl_151_n15), .B1(
        u1_adj_op_27_), .B2(u1_srl_151_n16), .ZN(u1_srl_151_n341) );
  OAI221_X1 u1_srl_151_U377 ( .B1(u1_srl_151_n7), .B2(u1_srl_151_n116), .C1(
        u1_srl_151_n12), .C2(u1_srl_151_n115), .A(u1_srl_151_n341), .ZN(
        u1_srl_151_n259) );
  AOI22_X1 u1_srl_151_U376 ( .A1(n6252), .A2(u1_srl_151_n15), .B1(n6255), .B2(
        u1_srl_151_n16), .ZN(u1_srl_151_n340) );
  OAI221_X1 u1_srl_151_U375 ( .B1(u1_srl_151_n7), .B2(u1_srl_151_n120), .C1(
        u1_srl_151_n12), .C2(u1_srl_151_n119), .A(u1_srl_151_n340), .ZN(
        u1_srl_151_n255) );
  AOI22_X1 u1_srl_151_U374 ( .A1(u1_adj_op_38_), .A2(u1_srl_151_n15), .B1(
        n6245), .B2(u1_srl_151_n16), .ZN(u1_srl_151_n339) );
  OAI221_X1 u1_srl_151_U373 ( .B1(u1_srl_151_n7), .B2(u1_srl_151_n107), .C1(
        u1_srl_151_n12), .C2(u1_srl_151_n106), .A(u1_srl_151_n339), .ZN(
        u1_srl_151_n260) );
  AOI22_X1 u1_srl_151_U372 ( .A1(n6246), .A2(u1_srl_151_n198), .B1(n6248), 
        .B2(u1_srl_151_n16), .ZN(u1_srl_151_n338) );
  OAI221_X1 u1_srl_151_U371 ( .B1(u1_srl_151_n7), .B2(u1_srl_151_n111), .C1(
        u1_srl_151_n12), .C2(u1_srl_151_n110), .A(u1_srl_151_n338), .ZN(
        u1_srl_151_n258) );
  AOI22_X1 u1_srl_151_U370 ( .A1(u1_srl_151_n237), .A2(u1_srl_151_n260), .B1(
        u1_srl_151_n196), .B2(u1_srl_151_n258), .ZN(u1_srl_151_n337) );
  AOI221_X1 u1_srl_151_U369 ( .B1(u1_srl_151_n259), .B2(u1_srl_151_n11), .C1(
        u1_srl_151_n255), .C2(u1_srl_151_n2), .A(u1_srl_151_n48), .ZN(
        u1_srl_151_n231) );
  AOI22_X1 u1_srl_151_U368 ( .A1(n6239), .A2(u1_srl_151_n15), .B1(n6241), .B2(
        u1_srl_151_n16), .ZN(u1_srl_151_n336) );
  AOI221_X1 u1_srl_151_U367 ( .B1(u1_srl_151_n224), .B2(u1_adj_op_44_), .C1(
        u1_srl_151_n13), .C2(n6240), .A(u1_srl_151_n69), .ZN(u1_srl_151_n263)
         );
  AOI22_X1 u1_srl_151_U366 ( .A1(u1_adj_op_42_), .A2(u1_srl_151_n15), .B1(
        n6244), .B2(u1_srl_151_n16), .ZN(u1_srl_151_n335) );
  AOI221_X1 u1_srl_151_U365 ( .B1(u1_srl_151_n224), .B2(n6243), .C1(
        u1_srl_151_n13), .C2(n6242), .A(u1_srl_151_n71), .ZN(u1_srl_151_n286)
         );
  AOI22_X1 u1_srl_151_U364 ( .A1(u1_srl_151_n16), .A2(u1_adj_op_51_), .B1(
        u1_srl_151_n224), .B2(n4266), .ZN(u1_srl_151_n177) );
  AOI22_X1 u1_srl_151_U363 ( .A1(n6234), .A2(u1_srl_151_n15), .B1(n6238), .B2(
        u1_srl_151_n16), .ZN(u1_srl_151_n334) );
  AOI221_X1 u1_srl_151_U362 ( .B1(u1_srl_151_n224), .B2(n6237), .C1(
        u1_srl_151_n13), .C2(n6236), .A(u1_srl_151_n74), .ZN(u1_srl_151_n262)
         );
  OAI22_X1 u1_srl_151_U361 ( .A1(u1_srl_151_n58), .A2(u1_srl_151_n177), .B1(
        u1_srl_151_n5), .B2(u1_srl_151_n262), .ZN(u1_srl_151_n333) );
  AOI221_X1 u1_srl_151_U360 ( .B1(u1_srl_151_n68), .B2(u1_srl_151_n11), .C1(
        u1_srl_151_n70), .C2(u1_srl_151_n2), .A(u1_srl_151_n333), .ZN(
        u1_srl_151_n191) );
  AOI22_X1 u1_srl_151_U359 ( .A1(u1_adj_op_10_), .A2(u1_srl_151_n198), .B1(
        n6231), .B2(u1_srl_151_n16), .ZN(u1_srl_151_n332) );
  OAI221_X1 u1_srl_151_U358 ( .B1(u1_srl_151_n7), .B2(u1_srl_151_n100), .C1(
        u1_srl_151_n12), .C2(u1_srl_151_n99), .A(u1_srl_151_n332), .ZN(
        u1_srl_151_n167) );
  AOI22_X1 u1_srl_151_U357 ( .A1(u1_srl_151_n145), .A2(u1_srl_151_n28), .B1(
        u1_srl_151_n146), .B2(u1_srl_151_n167), .ZN(u1_srl_151_n327) );
  AOI22_X1 u1_srl_151_U356 ( .A1(n6259), .A2(u1_srl_151_n198), .B1(
        u1_adj_op_11_), .B2(u1_srl_151_n16), .ZN(u1_srl_151_n331) );
  OAI221_X1 u1_srl_151_U355 ( .B1(u1_srl_151_n6), .B2(u1_srl_151_n133), .C1(
        u1_srl_151_n12), .C2(u1_srl_151_n132), .A(u1_srl_151_n331), .ZN(
        u1_srl_151_n169) );
  AOI22_X1 u1_srl_151_U354 ( .A1(u1_adj_op_22_), .A2(u1_srl_151_n198), .B1(
        u1_srl_151_n199), .B2(n6257), .ZN(u1_srl_151_n330) );
  OAI221_X1 u1_srl_151_U353 ( .B1(u1_srl_151_n6), .B2(u1_srl_151_n124), .C1(
        u1_srl_151_n12), .C2(u1_srl_151_n123), .A(u1_srl_151_n330), .ZN(
        u1_srl_151_n256) );
  AOI22_X1 u1_srl_151_U352 ( .A1(n6258), .A2(u1_srl_151_n198), .B1(
        u1_adj_op_15_), .B2(u1_srl_151_n16), .ZN(u1_srl_151_n329) );
  OAI221_X1 u1_srl_151_U351 ( .B1(u1_srl_151_n6), .B2(u1_srl_151_n129), .C1(
        u1_srl_151_n12), .C2(u1_srl_151_n128), .A(u1_srl_151_n329), .ZN(
        u1_srl_151_n168) );
  AOI222_X1 u1_srl_151_U350 ( .A1(u1_srl_151_n139), .A2(u1_srl_151_n169), .B1(
        u1_srl_151_n141), .B2(u1_srl_151_n256), .C1(u1_srl_151_n143), .C2(
        u1_srl_151_n168), .ZN(u1_srl_151_n328) );
  OAI211_X1 u1_srl_151_U349 ( .C1(u1_srl_151_n231), .C2(u1_srl_151_n96), .A(
        u1_srl_151_n327), .B(u1_srl_151_n328), .ZN(u1_adj_op_out_sft_10_) );
  AOI22_X1 u1_srl_151_U348 ( .A1(n6248), .A2(u1_srl_151_n198), .B1(
        u1_adj_op_28_), .B2(u1_srl_151_n16), .ZN(u1_srl_151_n326) );
  OAI221_X1 u1_srl_151_U347 ( .B1(u1_srl_151_n6), .B2(u1_srl_151_n115), .C1(
        u1_srl_151_n12), .C2(u1_srl_151_n113), .A(u1_srl_151_n326), .ZN(
        u1_srl_151_n279) );
  AOI22_X1 u1_srl_151_U346 ( .A1(u1_adj_op_27_), .A2(u1_srl_151_n15), .B1(
        n6254), .B2(u1_srl_151_n16), .ZN(u1_srl_151_n325) );
  OAI221_X1 u1_srl_151_U345 ( .B1(u1_srl_151_n6), .B2(u1_srl_151_n119), .C1(
        u1_srl_151_n12), .C2(u1_srl_151_n118), .A(u1_srl_151_n325), .ZN(
        u1_srl_151_n248) );
  AOI22_X1 u1_srl_151_U344 ( .A1(n6244), .A2(u1_srl_151_n15), .B1(
        u1_adj_op_36_), .B2(u1_srl_151_n16), .ZN(u1_srl_151_n324) );
  AOI221_X1 u1_srl_151_U343 ( .B1(u1_srl_151_n224), .B2(u1_adj_op_37_), .C1(
        u1_srl_151_n13), .C2(u1_adj_op_38_), .A(u1_srl_151_n78), .ZN(
        u1_srl_151_n283) );
  AOI22_X1 u1_srl_151_U342 ( .A1(n6245), .A2(u1_srl_151_n198), .B1(
        u1_adj_op_32_), .B2(u1_srl_151_n16), .ZN(u1_srl_151_n323) );
  OAI221_X1 u1_srl_151_U341 ( .B1(u1_srl_151_n6), .B2(u1_srl_151_n110), .C1(
        u1_srl_151_n12), .C2(u1_srl_151_n109), .A(u1_srl_151_n323), .ZN(
        u1_srl_151_n281) );
  OAI22_X1 u1_srl_151_U340 ( .A1(u1_srl_151_n58), .A2(u1_srl_151_n283), .B1(
        u1_srl_151_n5), .B2(u1_srl_151_n79), .ZN(u1_srl_151_n322) );
  AOI221_X1 u1_srl_151_U339 ( .B1(u1_srl_151_n279), .B2(u1_srl_151_n11), .C1(
        u1_srl_151_n248), .C2(u1_srl_151_n2), .A(u1_srl_151_n322), .ZN(
        u1_srl_151_n229) );
  AOI22_X1 u1_srl_151_U338 ( .A1(n6241), .A2(u1_srl_151_n15), .B1(n6243), .B2(
        u1_srl_151_n16), .ZN(u1_srl_151_n321) );
  AOI221_X1 u1_srl_151_U337 ( .B1(u1_srl_151_n224), .B2(n6242), .C1(
        u1_srl_151_n13), .C2(u1_adj_op_42_), .A(u1_srl_151_n81), .ZN(
        u1_srl_151_n254) );
  AOI22_X1 u1_srl_151_U336 ( .A1(n6238), .A2(u1_srl_151_n15), .B1(
        u1_adj_op_44_), .B2(u1_srl_151_n16), .ZN(u1_srl_151_n320) );
  AOI221_X1 u1_srl_151_U335 ( .B1(u1_srl_151_n224), .B2(n6240), .C1(
        u1_srl_151_n13), .C2(n6239), .A(u1_srl_151_n82), .ZN(u1_srl_151_n253)
         );
  NAND2_X1 u1_srl_151_U334 ( .A1(n4266), .A2(u1_srl_151_n199), .ZN(
        u1_srl_151_n176) );
  AOI22_X1 u1_srl_151_U333 ( .A1(u1_adj_op_51_), .A2(u1_srl_151_n15), .B1(
        n6237), .B2(u1_srl_151_n16), .ZN(u1_srl_151_n319) );
  AOI221_X1 u1_srl_151_U332 ( .B1(u1_srl_151_n224), .B2(n6236), .C1(
        u1_srl_151_n13), .C2(n6234), .A(u1_srl_151_n83), .ZN(u1_srl_151_n252)
         );
  MUX2_X1 u1_srl_151_U331 ( .A(u1_srl_151_n176), .B(u1_srl_151_n252), .S(
        u1_srl_151_n59), .Z(u1_srl_151_n280) );
  OAI222_X1 u1_srl_151_U330 ( .A1(u1_srl_151_n254), .A2(u1_srl_151_n19), .B1(
        u1_srl_151_n253), .B2(u1_srl_151_n1), .C1(u1_srl_151_n280), .C2(
        u1_srl_151_n94), .ZN(u1_srl_151_n230) );
  AOI22_X1 u1_srl_151_U329 ( .A1(u1_adj_op_11_), .A2(u1_srl_151_n15), .B1(
        n6230), .B2(u1_srl_151_n16), .ZN(u1_srl_151_n318) );
  OAI221_X1 u1_srl_151_U328 ( .B1(u1_srl_151_n6), .B2(u1_srl_151_n99), .C1(
        u1_srl_151_n12), .C2(u1_srl_151_n135), .A(u1_srl_151_n318), .ZN(
        u1_srl_151_n159) );
  AOI22_X1 u1_srl_151_U327 ( .A1(u1_srl_151_n145), .A2(u1_srl_151_n230), .B1(
        u1_srl_151_n146), .B2(u1_srl_151_n159), .ZN(u1_srl_151_n313) );
  AOI22_X1 u1_srl_151_U326 ( .A1(u1_adj_op_15_), .A2(u1_srl_151_n15), .B1(
        n6261), .B2(u1_srl_151_n16), .ZN(u1_srl_151_n317) );
  OAI221_X1 u1_srl_151_U325 ( .B1(u1_srl_151_n6), .B2(u1_srl_151_n132), .C1(
        u1_srl_151_n12), .C2(u1_srl_151_n131), .A(u1_srl_151_n317), .ZN(
        u1_srl_151_n161) );
  AOI22_X1 u1_srl_151_U324 ( .A1(n6255), .A2(u1_srl_151_n15), .B1(
        u1_srl_151_n199), .B2(u1_adj_op_20_), .ZN(u1_srl_151_n316) );
  OAI221_X1 u1_srl_151_U323 ( .B1(u1_srl_151_n6), .B2(u1_srl_151_n123), .C1(
        u1_srl_151_n12), .C2(u1_srl_151_n122), .A(u1_srl_151_n316), .ZN(
        u1_srl_151_n249) );
  AOI22_X1 u1_srl_151_U322 ( .A1(u1_srl_151_n15), .A2(n6257), .B1(
        u1_adj_op_16_), .B2(u1_srl_151_n16), .ZN(u1_srl_151_n315) );
  OAI221_X1 u1_srl_151_U321 ( .B1(u1_srl_151_n6), .B2(u1_srl_151_n128), .C1(
        u1_srl_151_n12), .C2(u1_srl_151_n127), .A(u1_srl_151_n315), .ZN(
        u1_srl_151_n160) );
  AOI222_X1 u1_srl_151_U320 ( .A1(u1_srl_151_n139), .A2(u1_srl_151_n161), .B1(
        u1_srl_151_n141), .B2(u1_srl_151_n249), .C1(u1_srl_151_n143), .C2(
        u1_srl_151_n160), .ZN(u1_srl_151_n314) );
  OAI211_X1 u1_srl_151_U319 ( .C1(u1_srl_151_n229), .C2(u1_srl_151_n96), .A(
        u1_srl_151_n313), .B(u1_srl_151_n314), .ZN(u1_adj_op_out_sft_11_) );
  AOI22_X1 u1_srl_151_U318 ( .A1(u1_srl_151_n237), .A2(u1_srl_151_n62), .B1(
        u1_srl_151_n196), .B2(u1_srl_151_n245), .ZN(u1_srl_151_n311) );
  AOI221_X1 u1_srl_151_U317 ( .B1(u1_srl_151_n246), .B2(u1_srl_151_n11), .C1(
        u1_srl_151_n242), .C2(u1_srl_151_n2), .A(u1_srl_151_n49), .ZN(
        u1_srl_151_n228) );
  AOI222_X1 u1_srl_151_U316 ( .A1(u1_srl_151_n64), .A2(u1_srl_151_n10), .B1(
        u1_srl_151_n66), .B2(u1_srl_151_n196), .C1(u1_srl_151_n60), .C2(
        u1_srl_151_n2), .ZN(u1_srl_151_n190) );
  AOI22_X1 u1_srl_151_U315 ( .A1(u1_srl_151_n145), .A2(u1_srl_151_n29), .B1(
        u1_srl_151_n146), .B2(u1_srl_151_n152), .ZN(u1_srl_151_n309) );
  AOI222_X1 u1_srl_151_U314 ( .A1(u1_srl_151_n139), .A2(u1_srl_151_n154), .B1(
        u1_srl_151_n141), .B2(u1_srl_151_n243), .C1(u1_srl_151_n143), .C2(
        u1_srl_151_n153), .ZN(u1_srl_151_n310) );
  OAI211_X1 u1_srl_151_U313 ( .C1(u1_srl_151_n228), .C2(u1_srl_151_n96), .A(
        u1_srl_151_n309), .B(u1_srl_151_n310), .ZN(u1_adj_op_out_sft_12_) );
  AOI22_X1 u1_srl_151_U312 ( .A1(n6247), .A2(u1_srl_151_n15), .B1(n6249), .B2(
        u1_srl_151_n16), .ZN(u1_srl_151_n308) );
  OAI221_X1 u1_srl_151_U311 ( .B1(u1_srl_151_n6), .B2(u1_srl_151_n112), .C1(
        u1_srl_151_n12), .C2(u1_srl_151_n111), .A(u1_srl_151_n308), .ZN(
        u1_srl_151_n239) );
  AOI22_X1 u1_srl_151_U310 ( .A1(n6251), .A2(u1_srl_151_n15), .B1(n6252), .B2(
        u1_srl_151_n16), .ZN(u1_srl_151_n307) );
  OAI221_X1 u1_srl_151_U309 ( .B1(u1_srl_151_n6), .B2(u1_srl_151_n117), .C1(
        u1_srl_151_n3), .C2(u1_srl_151_n116), .A(u1_srl_151_n307), .ZN(
        u1_srl_151_n234) );
  AOI22_X1 u1_srl_151_U308 ( .A1(n6242), .A2(u1_srl_151_n15), .B1(
        u1_adj_op_38_), .B2(u1_srl_151_n16), .ZN(u1_srl_151_n306) );
  AOI221_X1 u1_srl_151_U307 ( .B1(u1_srl_151_n224), .B2(n6244), .C1(
        u1_srl_151_n13), .C2(n6243), .A(u1_srl_151_n86), .ZN(u1_srl_151_n267)
         );
  AOI22_X1 u1_srl_151_U306 ( .A1(u1_adj_op_37_), .A2(u1_srl_151_n15), .B1(
        n6246), .B2(u1_srl_151_n16), .ZN(u1_srl_151_n305) );
  OAI221_X1 u1_srl_151_U305 ( .B1(u1_srl_151_n6), .B2(u1_srl_151_n108), .C1(
        u1_srl_151_n3), .C2(u1_srl_151_n107), .A(u1_srl_151_n305), .ZN(
        u1_srl_151_n238) );
  OAI22_X1 u1_srl_151_U304 ( .A1(u1_srl_151_n58), .A2(u1_srl_151_n267), .B1(
        u1_srl_151_n5), .B2(u1_srl_151_n87), .ZN(u1_srl_151_n304) );
  AOI221_X1 u1_srl_151_U303 ( .B1(u1_srl_151_n239), .B2(u1_srl_151_n11), .C1(
        u1_srl_151_n234), .C2(u1_srl_151_n2), .A(u1_srl_151_n304), .ZN(
        u1_srl_151_n227) );
  AOI22_X1 u1_srl_151_U302 ( .A1(n6236), .A2(u1_srl_151_n15), .B1(n6239), .B2(
        u1_srl_151_n16), .ZN(u1_srl_151_n303) );
  AOI221_X1 u1_srl_151_U301 ( .B1(u1_srl_151_n224), .B2(n6238), .C1(
        u1_srl_151_n13), .C2(n6237), .A(u1_srl_151_n89), .ZN(u1_srl_151_n233)
         );
  AOI222_X1 u1_srl_151_U300 ( .A1(u1_srl_151_n13), .A2(n4266), .B1(
        u1_srl_151_n224), .B2(u1_adj_op_51_), .C1(u1_srl_151_n16), .C2(n6234), 
        .ZN(u1_srl_151_n178) );
  AOI22_X1 u1_srl_151_U299 ( .A1(n6240), .A2(u1_srl_151_n15), .B1(
        u1_adj_op_42_), .B2(u1_srl_151_n16), .ZN(u1_srl_151_n302) );
  AOI221_X1 u1_srl_151_U298 ( .B1(u1_srl_151_n224), .B2(n6241), .C1(
        u1_srl_151_n13), .C2(u1_adj_op_44_), .A(u1_srl_151_n92), .ZN(
        u1_srl_151_n266) );
  AOI222_X1 u1_srl_151_U297 ( .A1(u1_srl_151_n88), .A2(u1_srl_151_n10), .B1(
        u1_srl_151_n90), .B2(u1_srl_151_n196), .C1(u1_srl_151_n91), .C2(
        u1_srl_151_n2), .ZN(u1_srl_151_n189) );
  AOI22_X1 u1_srl_151_U296 ( .A1(n6260), .A2(u1_srl_151_n15), .B1(
        u1_adj_op_10_), .B2(u1_srl_151_n199), .ZN(u1_srl_151_n301) );
  OAI221_X1 u1_srl_151_U295 ( .B1(u1_srl_151_n6), .B2(u1_srl_151_n134), .C1(
        u1_srl_151_n3), .C2(u1_srl_151_n133), .A(u1_srl_151_n301), .ZN(
        u1_srl_151_n140) );
  AOI22_X1 u1_srl_151_U294 ( .A1(u1_srl_151_n145), .A2(u1_srl_151_n30), .B1(
        u1_srl_151_n146), .B2(u1_srl_151_n140), .ZN(u1_srl_151_n296) );
  AOI22_X1 u1_srl_151_U293 ( .A1(u1_adj_op_17_), .A2(u1_srl_151_n15), .B1(
        n6259), .B2(u1_srl_151_n199), .ZN(u1_srl_151_n300) );
  OAI221_X1 u1_srl_151_U292 ( .B1(u1_srl_151_n6), .B2(u1_srl_151_n130), .C1(
        u1_srl_151_n3), .C2(u1_srl_151_n129), .A(u1_srl_151_n300), .ZN(
        u1_srl_151_n144) );
  AOI22_X1 u1_srl_151_U291 ( .A1(n6253), .A2(u1_srl_151_n15), .B1(
        u1_adj_op_22_), .B2(u1_srl_151_n16), .ZN(u1_srl_151_n299) );
  OAI221_X1 u1_srl_151_U290 ( .B1(u1_srl_151_n6), .B2(u1_srl_151_n121), .C1(
        u1_srl_151_n3), .C2(u1_srl_151_n120), .A(u1_srl_151_n299), .ZN(
        u1_srl_151_n235) );
  AOI22_X1 u1_srl_151_U289 ( .A1(u1_adj_op_21_), .A2(u1_srl_151_n15), .B1(
        n6258), .B2(u1_srl_151_n16), .ZN(u1_srl_151_n298) );
  OAI221_X1 u1_srl_151_U288 ( .B1(u1_srl_151_n6), .B2(u1_srl_151_n126), .C1(
        u1_srl_151_n3), .C2(u1_srl_151_n124), .A(u1_srl_151_n298), .ZN(
        u1_srl_151_n142) );
  AOI222_X1 u1_srl_151_U287 ( .A1(u1_srl_151_n139), .A2(u1_srl_151_n144), .B1(
        u1_srl_151_n141), .B2(u1_srl_151_n235), .C1(u1_srl_151_n143), .C2(
        u1_srl_151_n142), .ZN(u1_srl_151_n297) );
  OAI211_X1 u1_srl_151_U286 ( .C1(u1_srl_151_n227), .C2(u1_srl_151_n96), .A(
        u1_srl_151_n296), .B(u1_srl_151_n297), .ZN(u1_adj_op_out_sft_13_) );
  AOI22_X1 u1_srl_151_U285 ( .A1(u1_srl_151_n237), .A2(u1_srl_151_n70), .B1(
        u1_srl_151_n196), .B2(u1_srl_151_n260), .ZN(u1_srl_151_n295) );
  AOI221_X1 u1_srl_151_U284 ( .B1(u1_srl_151_n258), .B2(u1_srl_151_n10), .C1(
        u1_srl_151_n259), .C2(u1_srl_151_n18), .A(u1_srl_151_n50), .ZN(
        u1_srl_151_n218) );
  AOI222_X1 u1_srl_151_U283 ( .A1(u1_srl_151_n73), .A2(u1_srl_151_n10), .B1(
        u1_srl_151_n72), .B2(u1_srl_151_n196), .C1(u1_srl_151_n68), .C2(
        u1_srl_151_n2), .ZN(u1_srl_151_n188) );
  AOI22_X1 u1_srl_151_U282 ( .A1(u1_srl_151_n145), .A2(u1_srl_151_n31), .B1(
        u1_srl_151_n146), .B2(u1_srl_151_n169), .ZN(u1_srl_151_n293) );
  AOI222_X1 u1_srl_151_U281 ( .A1(u1_srl_151_n139), .A2(u1_srl_151_n168), .B1(
        u1_srl_151_n141), .B2(u1_srl_151_n255), .C1(u1_srl_151_n143), .C2(
        u1_srl_151_n256), .ZN(u1_srl_151_n294) );
  OAI211_X1 u1_srl_151_U280 ( .C1(u1_srl_151_n218), .C2(u1_srl_151_n96), .A(
        u1_srl_151_n293), .B(u1_srl_151_n294), .ZN(u1_adj_op_out_sft_14_) );
  OAI22_X1 u1_srl_151_U279 ( .A1(u1_srl_151_n58), .A2(u1_srl_151_n254), .B1(
        u1_srl_151_n5), .B2(u1_srl_151_n283), .ZN(u1_srl_151_n292) );
  AOI221_X1 u1_srl_151_U278 ( .B1(u1_srl_151_n281), .B2(u1_srl_151_n11), .C1(
        u1_srl_151_n279), .C2(u1_srl_151_n2), .A(u1_srl_151_n292), .ZN(
        u1_srl_151_n216) );
  OAI222_X1 u1_srl_151_U277 ( .A1(u1_srl_151_n252), .A2(u1_srl_151_n1), .B1(
        u1_srl_151_n5), .B2(u1_srl_151_n176), .C1(u1_srl_151_n253), .C2(
        u1_srl_151_n19), .ZN(u1_srl_151_n217) );
  AOI22_X1 u1_srl_151_U276 ( .A1(u1_srl_151_n145), .A2(u1_srl_151_n217), .B1(
        u1_srl_151_n146), .B2(u1_srl_151_n161), .ZN(u1_srl_151_n290) );
  AOI222_X1 u1_srl_151_U275 ( .A1(u1_srl_151_n139), .A2(u1_srl_151_n160), .B1(
        u1_srl_151_n141), .B2(u1_srl_151_n248), .C1(u1_srl_151_n143), .C2(
        u1_srl_151_n249), .ZN(u1_srl_151_n291) );
  OAI211_X1 u1_srl_151_U274 ( .C1(u1_srl_151_n216), .C2(u1_srl_151_n96), .A(
        u1_srl_151_n290), .B(u1_srl_151_n291), .ZN(u1_adj_op_out_sft_15_) );
  OAI222_X1 u1_srl_151_U273 ( .A1(u1_srl_151_n215), .A2(u1_srl_151_n96), .B1(
        u1_srl_151_n187), .B2(u1_srl_151_n95), .C1(u1_srl_151_n289), .C2(
        u1_srl_151_n9), .ZN(u1_adj_op_out_sft_16_) );
  OAI22_X1 u1_srl_151_U272 ( .A1(u1_srl_151_n58), .A2(u1_srl_151_n266), .B1(
        u1_srl_151_n5), .B2(u1_srl_151_n267), .ZN(u1_srl_151_n288) );
  AOI221_X1 u1_srl_151_U271 ( .B1(u1_srl_151_n238), .B2(u1_srl_151_n11), .C1(
        u1_srl_151_n239), .C2(u1_srl_151_n18), .A(u1_srl_151_n288), .ZN(
        u1_srl_151_n214) );
  AOI22_X1 u1_srl_151_U270 ( .A1(u1_srl_151_n88), .A2(u1_srl_151_n2), .B1(
        u1_srl_151_n90), .B2(u1_srl_151_n11), .ZN(u1_srl_151_n186) );
  AOI22_X1 u1_srl_151_U269 ( .A1(u1_srl_151_n237), .A2(u1_srl_151_n234), .B1(
        u1_srl_151_n196), .B2(u1_srl_151_n235), .ZN(u1_srl_151_n287) );
  AOI221_X1 u1_srl_151_U268 ( .B1(u1_srl_151_n142), .B2(u1_srl_151_n10), .C1(
        u1_srl_151_n144), .C2(u1_srl_151_n18), .A(u1_srl_151_n51), .ZN(
        u1_srl_151_n277) );
  OAI222_X1 u1_srl_151_U267 ( .A1(u1_srl_151_n214), .A2(u1_srl_151_n96), .B1(
        u1_srl_151_n186), .B2(u1_srl_151_n95), .C1(u1_srl_151_n277), .C2(
        u1_srl_151_n9), .ZN(u1_adj_op_out_sft_17_) );
  OAI22_X1 u1_srl_151_U266 ( .A1(u1_srl_151_n58), .A2(u1_srl_151_n263), .B1(
        u1_srl_151_n5), .B2(u1_srl_151_n286), .ZN(u1_srl_151_n285) );
  AOI221_X1 u1_srl_151_U265 ( .B1(u1_srl_151_n260), .B2(u1_srl_151_n10), .C1(
        u1_srl_151_n258), .C2(u1_srl_151_n18), .A(u1_srl_151_n285), .ZN(
        u1_srl_151_n213) );
  AOI22_X1 u1_srl_151_U264 ( .A1(u1_srl_151_n73), .A2(u1_srl_151_n18), .B1(
        u1_srl_151_n72), .B2(u1_srl_151_n11), .ZN(u1_srl_151_n181) );
  AOI22_X1 u1_srl_151_U263 ( .A1(u1_srl_151_n237), .A2(u1_srl_151_n259), .B1(
        u1_srl_151_n196), .B2(u1_srl_151_n255), .ZN(u1_srl_151_n284) );
  AOI221_X1 u1_srl_151_U262 ( .B1(u1_srl_151_n256), .B2(u1_srl_151_n10), .C1(
        u1_srl_151_n168), .C2(u1_srl_151_n18), .A(u1_srl_151_n52), .ZN(
        u1_srl_151_n226) );
  OAI222_X1 u1_srl_151_U261 ( .A1(u1_srl_151_n213), .A2(u1_srl_151_n96), .B1(
        u1_srl_151_n181), .B2(u1_srl_151_n95), .C1(u1_srl_151_n226), .C2(
        u1_srl_151_n9), .ZN(u1_adj_op_out_sft_18_) );
  OAI22_X1 u1_srl_151_U260 ( .A1(u1_srl_151_n58), .A2(u1_srl_151_n253), .B1(
        u1_srl_151_n5), .B2(u1_srl_151_n254), .ZN(u1_srl_151_n282) );
  AOI221_X1 u1_srl_151_U259 ( .B1(u1_srl_151_n77), .B2(u1_srl_151_n11), .C1(
        u1_srl_151_n281), .C2(u1_srl_151_n18), .A(u1_srl_151_n282), .ZN(
        u1_srl_151_n212) );
  OR2_X1 u1_srl_151_U258 ( .A1(u1_srl_151_n280), .A2(n6224), .ZN(
        u1_srl_151_n180) );
  OAI22_X1 u1_srl_151_U257 ( .A1(u1_srl_151_n58), .A2(u1_srl_151_n75), .B1(
        u1_srl_151_n5), .B2(u1_srl_151_n76), .ZN(u1_srl_151_n278) );
  AOI221_X1 u1_srl_151_U256 ( .B1(u1_srl_151_n249), .B2(u1_srl_151_n10), .C1(
        u1_srl_151_n160), .C2(u1_srl_151_n18), .A(u1_srl_151_n278), .ZN(
        u1_srl_151_n201) );
  OAI222_X1 u1_srl_151_U255 ( .A1(u1_srl_151_n212), .A2(u1_srl_151_n96), .B1(
        u1_srl_151_n95), .B2(u1_srl_151_n180), .C1(u1_srl_151_n201), .C2(
        u1_srl_151_n9), .ZN(u1_adj_op_out_sft_19_) );
  AOI22_X1 u1_srl_151_U254 ( .A1(n6233), .A2(u1_srl_151_n15), .B1(n6250), .B2(
        u1_srl_151_n199), .ZN(u1_srl_151_n276) );
  OAI221_X1 u1_srl_151_U253 ( .B1(u1_srl_151_n6), .B2(u1_srl_151_n105), .C1(
        u1_srl_151_n3), .C2(u1_srl_151_n104), .A(u1_srl_151_n276), .ZN(
        u1_srl_151_n174) );
  AOI222_X1 u1_srl_151_U252 ( .A1(u1_srl_151_n163), .A2(u1_srl_151_n33), .B1(
        u1_srl_151_n139), .B2(u1_srl_151_n174), .C1(u1_srl_151_n145), .C2(
        u1_srl_151_n32), .ZN(u1_srl_151_n271) );
  AOI22_X1 u1_srl_151_U251 ( .A1(u1_srl_151_n15), .A2(n6256), .B1(
        u1_srl_151_n13), .B2(u1_adj_op_0_), .ZN(u1_srl_151_n273) );
  AOI22_X1 u1_srl_151_U250 ( .A1(n6229), .A2(u1_srl_151_n15), .B1(n6232), .B2(
        u1_srl_151_n199), .ZN(u1_srl_151_n275) );
  OAI221_X1 u1_srl_151_U249 ( .B1(u1_srl_151_n6), .B2(u1_srl_151_n101), .C1(
        u1_srl_151_n3), .C2(u1_srl_151_n100), .A(u1_srl_151_n275), .ZN(
        u1_srl_151_n147) );
  AOI22_X1 u1_srl_151_U248 ( .A1(u1_srl_151_n147), .A2(u1_srl_151_n143), .B1(
        u1_srl_151_n140), .B2(u1_srl_151_n141), .ZN(u1_srl_151_n274) );
  OAI221_X1 u1_srl_151_U247 ( .B1(u1_srl_151_n25), .B2(u1_srl_151_n273), .C1(
        u1_srl_151_n223), .C2(u1_srl_151_n186), .A(u1_srl_151_n274), .ZN(
        u1_srl_151_n272) );
  NAND2_X1 u1_srl_151_U246 ( .A1(u1_srl_151_n271), .A2(u1_srl_151_n24), .ZN(
        u1_adj_op_out_sft_1_) );
  OAI22_X1 u1_srl_151_U245 ( .A1(u1_srl_151_n58), .A2(u1_srl_151_n241), .B1(
        u1_srl_151_n5), .B2(u1_srl_151_n270), .ZN(u1_srl_151_n269) );
  AOI221_X1 u1_srl_151_U244 ( .B1(u1_srl_151_n62), .B2(u1_srl_151_n11), .C1(
        u1_srl_151_n245), .C2(u1_srl_151_n18), .A(u1_srl_151_n269), .ZN(
        u1_srl_151_n211) );
  NAND2_X1 u1_srl_151_U243 ( .A1(u1_srl_151_n145), .A2(u1_srl_151_n2), .ZN(
        u1_srl_151_n247) );
  AOI22_X1 u1_srl_151_U242 ( .A1(u1_srl_151_n237), .A2(u1_srl_151_n246), .B1(
        u1_srl_151_n196), .B2(u1_srl_151_n242), .ZN(u1_srl_151_n268) );
  AOI221_X1 u1_srl_151_U241 ( .B1(u1_srl_151_n243), .B2(u1_srl_151_n10), .C1(
        u1_srl_151_n153), .C2(u1_srl_151_n18), .A(u1_srl_151_n53), .ZN(
        u1_srl_151_n185) );
  OAI222_X1 u1_srl_151_U240 ( .A1(u1_srl_151_n211), .A2(u1_srl_151_n96), .B1(
        u1_srl_151_n179), .B2(u1_srl_151_n247), .C1(u1_srl_151_n185), .C2(
        u1_srl_151_n9), .ZN(u1_adj_op_out_sft_20_) );
  OAI22_X1 u1_srl_151_U239 ( .A1(u1_srl_151_n58), .A2(u1_srl_151_n233), .B1(
        u1_srl_151_n5), .B2(u1_srl_151_n266), .ZN(u1_srl_151_n265) );
  AOI221_X1 u1_srl_151_U238 ( .B1(u1_srl_151_n85), .B2(u1_srl_151_n11), .C1(
        u1_srl_151_n238), .C2(u1_srl_151_n18), .A(u1_srl_151_n265), .ZN(
        u1_srl_151_n209) );
  AOI22_X1 u1_srl_151_U237 ( .A1(u1_srl_151_n237), .A2(u1_srl_151_n239), .B1(
        u1_srl_151_n196), .B2(u1_srl_151_n234), .ZN(u1_srl_151_n264) );
  AOI221_X1 u1_srl_151_U236 ( .B1(u1_srl_151_n235), .B2(u1_srl_151_n10), .C1(
        u1_srl_151_n142), .C2(u1_srl_151_n2), .A(u1_srl_151_n54), .ZN(
        u1_srl_151_n175) );
  OAI222_X1 u1_srl_151_U235 ( .A1(u1_srl_151_n209), .A2(u1_srl_151_n96), .B1(
        u1_srl_151_n178), .B2(u1_srl_151_n247), .C1(u1_srl_151_n175), .C2(
        u1_srl_151_n9), .ZN(u1_adj_op_out_sft_21_) );
  OAI22_X1 u1_srl_151_U234 ( .A1(u1_srl_151_n58), .A2(u1_srl_151_n262), .B1(
        u1_srl_151_n5), .B2(u1_srl_151_n263), .ZN(u1_srl_151_n261) );
  AOI221_X1 u1_srl_151_U233 ( .B1(u1_srl_151_n70), .B2(u1_srl_151_n10), .C1(
        u1_srl_151_n260), .C2(u1_srl_151_n18), .A(u1_srl_151_n261), .ZN(
        u1_srl_151_n207) );
  AOI22_X1 u1_srl_151_U232 ( .A1(u1_srl_151_n237), .A2(u1_srl_151_n258), .B1(
        u1_srl_151_n196), .B2(u1_srl_151_n259), .ZN(u1_srl_151_n257) );
  AOI221_X1 u1_srl_151_U231 ( .B1(u1_srl_151_n255), .B2(u1_srl_151_n10), .C1(
        u1_srl_151_n256), .C2(u1_srl_151_n2), .A(u1_srl_151_n55), .ZN(
        u1_srl_151_n171) );
  OAI222_X1 u1_srl_151_U230 ( .A1(u1_srl_151_n207), .A2(u1_srl_151_n96), .B1(
        u1_srl_151_n177), .B2(u1_srl_151_n247), .C1(u1_srl_151_n171), .C2(
        u1_srl_151_n9), .ZN(u1_adj_op_out_sft_22_) );
  OAI22_X1 u1_srl_151_U229 ( .A1(u1_srl_151_n58), .A2(u1_srl_151_n252), .B1(
        u1_srl_151_n5), .B2(u1_srl_151_n253), .ZN(u1_srl_151_n251) );
  AOI221_X1 u1_srl_151_U228 ( .B1(u1_srl_151_n80), .B2(u1_srl_151_n10), .C1(
        u1_srl_151_n77), .C2(u1_srl_151_n2), .A(u1_srl_151_n251), .ZN(
        u1_srl_151_n204) );
  OAI22_X1 u1_srl_151_U227 ( .A1(u1_srl_151_n58), .A2(u1_srl_151_n79), .B1(
        u1_srl_151_n5), .B2(u1_srl_151_n75), .ZN(u1_srl_151_n250) );
  AOI221_X1 u1_srl_151_U226 ( .B1(u1_srl_151_n248), .B2(u1_srl_151_n10), .C1(
        u1_srl_151_n249), .C2(u1_srl_151_n2), .A(u1_srl_151_n250), .ZN(
        u1_srl_151_n164) );
  OAI222_X1 u1_srl_151_U225 ( .A1(u1_srl_151_n204), .A2(u1_srl_151_n96), .B1(
        u1_srl_151_n176), .B2(u1_srl_151_n247), .C1(u1_srl_151_n164), .C2(
        u1_srl_151_n9), .ZN(u1_adj_op_out_sft_23_) );
  AOI22_X1 u1_srl_151_U224 ( .A1(u1_srl_151_n237), .A2(u1_srl_151_n245), .B1(
        u1_srl_151_n196), .B2(u1_srl_151_n246), .ZN(u1_srl_151_n244) );
  AOI221_X1 u1_srl_151_U223 ( .B1(u1_srl_151_n242), .B2(u1_srl_151_n10), .C1(
        u1_srl_151_n243), .C2(u1_srl_151_n2), .A(u1_srl_151_n56), .ZN(
        u1_srl_151_n149) );
  OAI22_X1 u1_srl_151_U222 ( .A1(u1_srl_151_n58), .A2(u1_srl_151_n179), .B1(
        u1_srl_151_n5), .B2(u1_srl_151_n241), .ZN(u1_srl_151_n240) );
  AOI221_X1 u1_srl_151_U221 ( .B1(u1_srl_151_n60), .B2(u1_srl_151_n10), .C1(
        u1_srl_151_n62), .C2(u1_srl_151_n2), .A(u1_srl_151_n240), .ZN(
        u1_srl_151_n156) );
  OAI22_X1 u1_srl_151_U220 ( .A1(u1_srl_151_n149), .A2(u1_srl_151_n8), .B1(
        u1_srl_151_n156), .B2(u1_srl_151_n96), .ZN(u1_adj_op_out_sft_24_) );
  AOI22_X1 u1_srl_151_U219 ( .A1(u1_srl_151_n237), .A2(u1_srl_151_n238), .B1(
        u1_srl_151_n196), .B2(u1_srl_151_n239), .ZN(u1_srl_151_n236) );
  AOI221_X1 u1_srl_151_U218 ( .B1(u1_srl_151_n234), .B2(u1_srl_151_n10), .C1(
        u1_srl_151_n235), .C2(u1_srl_151_n2), .A(u1_srl_151_n57), .ZN(
        u1_srl_151_n136) );
  OAI22_X1 u1_srl_151_U217 ( .A1(u1_srl_151_n58), .A2(u1_srl_151_n178), .B1(
        u1_srl_151_n5), .B2(u1_srl_151_n233), .ZN(u1_srl_151_n232) );
  AOI221_X1 u1_srl_151_U216 ( .B1(u1_srl_151_n91), .B2(u1_srl_151_n10), .C1(
        u1_srl_151_n85), .C2(u1_srl_151_n2), .A(u1_srl_151_n232), .ZN(
        u1_srl_151_n148) );
  OAI22_X1 u1_srl_151_U215 ( .A1(u1_srl_151_n136), .A2(u1_srl_151_n8), .B1(
        u1_srl_151_n148), .B2(u1_srl_151_n96), .ZN(u1_adj_op_out_sft_25_) );
  OAI22_X1 u1_srl_151_U214 ( .A1(u1_srl_151_n231), .A2(u1_srl_151_n8), .B1(
        u1_srl_151_n191), .B2(u1_srl_151_n96), .ZN(u1_adj_op_out_sft_26_) );
  OAI22_X1 u1_srl_151_U213 ( .A1(u1_srl_151_n229), .A2(u1_srl_151_n8), .B1(
        u1_srl_151_n26), .B2(u1_srl_151_n96), .ZN(u1_adj_op_out_sft_27_) );
  OAI22_X1 u1_srl_151_U212 ( .A1(u1_srl_151_n228), .A2(u1_srl_151_n8), .B1(
        u1_srl_151_n190), .B2(u1_srl_151_n96), .ZN(u1_adj_op_out_sft_28_) );
  OAI22_X1 u1_srl_151_U211 ( .A1(u1_srl_151_n227), .A2(u1_srl_151_n8), .B1(
        u1_srl_151_n189), .B2(u1_srl_151_n96), .ZN(u1_adj_op_out_sft_29_) );
  AOI22_X1 u1_srl_151_U210 ( .A1(n6232), .A2(u1_srl_151_n15), .B1(u1_adj_op_3_), .B2(u1_srl_151_n199), .ZN(u1_srl_151_n225) );
  OAI221_X1 u1_srl_151_U209 ( .B1(u1_srl_151_n6), .B2(u1_srl_151_n104), .C1(
        u1_srl_151_n3), .C2(u1_srl_151_n103), .A(u1_srl_151_n225), .ZN(
        u1_srl_151_n170) );
  AOI222_X1 u1_srl_151_U208 ( .A1(u1_srl_151_n163), .A2(u1_srl_151_n35), .B1(
        u1_srl_151_n139), .B2(u1_srl_151_n170), .C1(u1_srl_151_n145), .C2(
        u1_srl_151_n34), .ZN(u1_srl_151_n219) );
  AOI222_X1 u1_srl_151_U207 ( .A1(n6250), .A2(u1_srl_151_n15), .B1(
        u1_adj_op_0_), .B2(u1_srl_151_n224), .C1(n6256), .C2(u1_srl_151_n13), 
        .ZN(u1_srl_151_n222) );
  OAI22_X1 u1_srl_151_U206 ( .A1(u1_srl_151_n222), .A2(u1_srl_151_n25), .B1(
        u1_srl_151_n181), .B2(u1_srl_151_n223), .ZN(u1_srl_151_n221) );
  AOI221_X1 u1_srl_151_U205 ( .B1(u1_srl_151_n141), .B2(u1_srl_151_n169), .C1(
        u1_srl_151_n143), .C2(u1_srl_151_n167), .A(u1_srl_151_n221), .ZN(
        u1_srl_151_n220) );
  NAND2_X1 u1_srl_151_U204 ( .A1(u1_srl_151_n219), .A2(u1_srl_151_n220), .ZN(
        u1_adj_op_out_sft_2_) );
  OAI22_X1 u1_srl_151_U203 ( .A1(u1_srl_151_n218), .A2(u1_srl_151_n8), .B1(
        u1_srl_151_n188), .B2(u1_srl_151_n96), .ZN(u1_adj_op_out_sft_30_) );
  OAI22_X1 u1_srl_151_U202 ( .A1(u1_srl_151_n216), .A2(u1_srl_151_n9), .B1(
        u1_srl_151_n27), .B2(u1_srl_151_n96), .ZN(u1_adj_op_out_sft_31_) );
  OAI22_X1 u1_srl_151_U201 ( .A1(u1_srl_151_n215), .A2(u1_srl_151_n8), .B1(
        u1_srl_151_n187), .B2(u1_srl_151_n96), .ZN(u1_adj_op_out_sft_32_) );
  OAI22_X1 u1_srl_151_U200 ( .A1(u1_srl_151_n214), .A2(u1_srl_151_n9), .B1(
        u1_srl_151_n186), .B2(u1_srl_151_n96), .ZN(u1_adj_op_out_sft_33_) );
  OAI22_X1 u1_srl_151_U199 ( .A1(u1_srl_151_n213), .A2(u1_srl_151_n9), .B1(
        u1_srl_151_n181), .B2(u1_srl_151_n96), .ZN(u1_adj_op_out_sft_34_) );
  MUX2_X1 u1_srl_151_U198 ( .A(u1_srl_151_n180), .B(u1_srl_151_n212), .S(
        u1_srl_151_n97), .Z(u1_srl_151_n202) );
  NOR2_X1 u1_srl_151_U197 ( .A1(n6226), .A2(u1_srl_151_n202), .ZN(
        u1_adj_op_out_sft_35_) );
  NAND2_X1 u1_srl_151_U196 ( .A1(n6225), .A2(u1_srl_151_n2), .ZN(
        u1_srl_151_n205) );
  OAI22_X1 u1_srl_151_U195 ( .A1(n6225), .A2(u1_srl_151_n211), .B1(
        u1_srl_151_n179), .B2(u1_srl_151_n205), .ZN(u1_srl_151_n210) );
  NOR2_X1 u1_srl_151_U194 ( .A1(n6226), .A2(u1_srl_151_n38), .ZN(
        u1_adj_op_out_sft_36_) );
  OAI22_X1 u1_srl_151_U193 ( .A1(n6225), .A2(u1_srl_151_n209), .B1(
        u1_srl_151_n178), .B2(u1_srl_151_n205), .ZN(u1_srl_151_n208) );
  NOR2_X1 u1_srl_151_U192 ( .A1(n6226), .A2(u1_srl_151_n40), .ZN(
        u1_adj_op_out_sft_37_) );
  OAI22_X1 u1_srl_151_U191 ( .A1(n6225), .A2(u1_srl_151_n207), .B1(
        u1_srl_151_n177), .B2(u1_srl_151_n205), .ZN(u1_srl_151_n206) );
  NOR2_X1 u1_srl_151_U190 ( .A1(n6226), .A2(u1_srl_151_n42), .ZN(
        u1_adj_op_out_sft_38_) );
  OAI22_X1 u1_srl_151_U189 ( .A1(n6225), .A2(u1_srl_151_n204), .B1(
        u1_srl_151_n205), .B2(u1_srl_151_n176), .ZN(u1_srl_151_n203) );
  NOR2_X1 u1_srl_151_U188 ( .A1(n6226), .A2(u1_srl_151_n44), .ZN(
        u1_adj_op_out_sft_39_) );
  OAI22_X1 u1_srl_151_U187 ( .A1(u1_srl_151_n3), .A2(u1_srl_151_n114), .B1(
        u1_srl_151_n6), .B2(u1_srl_151_n125), .ZN(u1_srl_151_n200) );
  AOI221_X1 u1_srl_151_U186 ( .B1(u1_adj_op_3_), .B2(u1_srl_151_n15), .C1(
        u1_adj_op_0_), .C2(u1_srl_151_n199), .A(u1_srl_151_n200), .ZN(
        u1_srl_151_n194) );
  AOI22_X1 u1_srl_151_U185 ( .A1(n6231), .A2(u1_srl_151_n198), .B1(n6235), 
        .B2(u1_srl_151_n16), .ZN(u1_srl_151_n197) );
  OAI221_X1 u1_srl_151_U184 ( .B1(u1_srl_151_n6), .B2(u1_srl_151_n103), .C1(
        u1_srl_151_n12), .C2(u1_srl_151_n102), .A(u1_srl_151_n197), .ZN(
        u1_srl_151_n162) );
  AOI22_X1 u1_srl_151_U183 ( .A1(u1_srl_151_n196), .A2(u1_srl_151_n159), .B1(
        u1_srl_151_n11), .B2(u1_srl_151_n162), .ZN(u1_srl_151_n195) );
  OAI221_X1 u1_srl_151_U182 ( .B1(u1_srl_151_n194), .B2(u1_srl_151_n19), .C1(
        u1_srl_151_n84), .C2(u1_srl_151_n58), .A(u1_srl_151_n195), .ZN(
        u1_srl_151_n193) );
  MUX2_X1 u1_srl_151_U181 ( .A(u1_srl_151_n37), .B(u1_srl_151_n193), .S(
        u1_srl_151_n97), .Z(u1_srl_151_n192) );
  MUX2_X1 u1_srl_151_U180 ( .A(u1_srl_151_n36), .B(u1_srl_151_n192), .S(
        u1_srl_151_n98), .Z(u1_adj_op_out_sft_3_) );
  NOR2_X1 u1_srl_151_U179 ( .A1(u1_srl_151_n156), .A2(u1_srl_151_n8), .ZN(
        u1_adj_op_out_sft_40_) );
  NOR2_X1 u1_srl_151_U178 ( .A1(u1_srl_151_n148), .A2(u1_srl_151_n8), .ZN(
        u1_adj_op_out_sft_41_) );
  NOR2_X1 u1_srl_151_U177 ( .A1(u1_srl_151_n191), .A2(u1_srl_151_n8), .ZN(
        u1_adj_op_out_sft_42_) );
  NOR2_X1 u1_srl_151_U176 ( .A1(u1_srl_151_n26), .A2(u1_srl_151_n8), .ZN(
        u1_adj_op_out_sft_43_) );
  NOR2_X1 u1_srl_151_U175 ( .A1(u1_srl_151_n190), .A2(u1_srl_151_n8), .ZN(
        u1_adj_op_out_sft_44_) );
  NOR2_X1 u1_srl_151_U174 ( .A1(u1_srl_151_n189), .A2(u1_srl_151_n8), .ZN(
        u1_adj_op_out_sft_45_) );
  NOR2_X1 u1_srl_151_U173 ( .A1(u1_srl_151_n188), .A2(u1_srl_151_n8), .ZN(
        u1_adj_op_out_sft_46_) );
  NOR2_X1 u1_srl_151_U172 ( .A1(u1_srl_151_n27), .A2(u1_srl_151_n8), .ZN(
        u1_adj_op_out_sft_47_) );
  NOR2_X1 u1_srl_151_U171 ( .A1(u1_srl_151_n187), .A2(u1_srl_151_n8), .ZN(
        u1_adj_op_out_sft_48_) );
  NOR2_X1 u1_srl_151_U170 ( .A1(u1_srl_151_n186), .A2(u1_srl_151_n8), .ZN(
        u1_adj_op_out_sft_49_) );
  AOI22_X1 u1_srl_151_U169 ( .A1(u1_srl_151_n146), .A2(u1_srl_151_n184), .B1(
        u1_srl_151_n163), .B2(u1_srl_151_n39), .ZN(u1_srl_151_n182) );
  AOI222_X1 u1_srl_151_U168 ( .A1(u1_srl_151_n139), .A2(u1_srl_151_n155), .B1(
        u1_srl_151_n141), .B2(u1_srl_151_n154), .C1(u1_srl_151_n143), .C2(
        u1_srl_151_n152), .ZN(u1_srl_151_n183) );
  OAI211_X1 u1_srl_151_U167 ( .C1(u1_srl_151_n38), .C2(u1_srl_151_n98), .A(
        u1_srl_151_n182), .B(u1_srl_151_n183), .ZN(u1_adj_op_out_sft_4_) );
  NOR2_X1 u1_srl_151_U166 ( .A1(u1_srl_151_n181), .A2(u1_srl_151_n8), .ZN(
        u1_adj_op_out_sft_50_) );
  NOR2_X1 u1_srl_151_U165 ( .A1(u1_srl_151_n8), .A2(u1_srl_151_n180), .ZN(
        u1_adj_op_out_sft_51_) );
  NOR2_X1 u1_srl_151_U164 ( .A1(u1_srl_151_n179), .A2(u1_srl_151_n25), .ZN(
        u1_adj_op_out_sft_52_) );
  NOR2_X1 u1_srl_151_U163 ( .A1(u1_srl_151_n178), .A2(u1_srl_151_n25), .ZN(
        u1_adj_op_out_sft_53_) );
  NOR2_X1 u1_srl_151_U162 ( .A1(u1_srl_151_n177), .A2(u1_srl_151_n25), .ZN(
        u1_adj_op_out_sft_54_) );
  NOR2_X1 u1_srl_151_U161 ( .A1(u1_srl_151_n25), .A2(u1_srl_151_n176), .ZN(
        u1_adj_op_out_sft_55_) );
  AOI22_X1 u1_srl_151_U160 ( .A1(u1_srl_151_n146), .A2(u1_srl_151_n174), .B1(
        u1_srl_151_n163), .B2(u1_srl_151_n41), .ZN(u1_srl_151_n172) );
  AOI222_X1 u1_srl_151_U159 ( .A1(u1_srl_151_n139), .A2(u1_srl_151_n147), .B1(
        u1_srl_151_n141), .B2(u1_srl_151_n144), .C1(u1_srl_151_n143), .C2(
        u1_srl_151_n140), .ZN(u1_srl_151_n173) );
  OAI211_X1 u1_srl_151_U158 ( .C1(u1_srl_151_n40), .C2(u1_srl_151_n98), .A(
        u1_srl_151_n172), .B(u1_srl_151_n173), .ZN(u1_adj_op_out_sft_5_) );
  AOI22_X1 u1_srl_151_U157 ( .A1(u1_srl_151_n146), .A2(u1_srl_151_n170), .B1(
        u1_srl_151_n163), .B2(u1_srl_151_n43), .ZN(u1_srl_151_n165) );
  AOI222_X1 u1_srl_151_U156 ( .A1(u1_srl_151_n139), .A2(u1_srl_151_n167), .B1(
        u1_srl_151_n141), .B2(u1_srl_151_n168), .C1(u1_srl_151_n143), .C2(
        u1_srl_151_n169), .ZN(u1_srl_151_n166) );
  OAI211_X1 u1_srl_151_U155 ( .C1(u1_srl_151_n42), .C2(u1_srl_151_n98), .A(
        u1_srl_151_n165), .B(u1_srl_151_n166), .ZN(u1_adj_op_out_sft_6_) );
  AOI22_X1 u1_srl_151_U154 ( .A1(u1_srl_151_n146), .A2(u1_srl_151_n162), .B1(
        u1_srl_151_n163), .B2(u1_srl_151_n45), .ZN(u1_srl_151_n157) );
  AOI222_X1 u1_srl_151_U153 ( .A1(u1_srl_151_n139), .A2(u1_srl_151_n159), .B1(
        u1_srl_151_n141), .B2(u1_srl_151_n160), .C1(u1_srl_151_n143), .C2(
        u1_srl_151_n161), .ZN(u1_srl_151_n158) );
  OAI211_X1 u1_srl_151_U152 ( .C1(u1_srl_151_n44), .C2(u1_srl_151_n98), .A(
        u1_srl_151_n157), .B(u1_srl_151_n158), .ZN(u1_adj_op_out_sft_7_) );
  AOI22_X1 u1_srl_151_U151 ( .A1(u1_srl_151_n145), .A2(u1_srl_151_n46), .B1(
        u1_srl_151_n146), .B2(u1_srl_151_n155), .ZN(u1_srl_151_n150) );
  AOI222_X1 u1_srl_151_U150 ( .A1(u1_srl_151_n139), .A2(u1_srl_151_n152), .B1(
        u1_srl_151_n141), .B2(u1_srl_151_n153), .C1(u1_srl_151_n143), .C2(
        u1_srl_151_n154), .ZN(u1_srl_151_n151) );
  OAI211_X1 u1_srl_151_U149 ( .C1(u1_srl_151_n149), .C2(u1_srl_151_n96), .A(
        u1_srl_151_n150), .B(u1_srl_151_n151), .ZN(u1_adj_op_out_sft_8_) );
  AOI22_X1 u1_srl_151_U148 ( .A1(u1_srl_151_n145), .A2(u1_srl_151_n47), .B1(
        u1_srl_151_n146), .B2(u1_srl_151_n147), .ZN(u1_srl_151_n137) );
  AOI222_X1 u1_srl_151_U147 ( .A1(u1_srl_151_n139), .A2(u1_srl_151_n140), .B1(
        u1_srl_151_n141), .B2(u1_srl_151_n142), .C1(u1_srl_151_n143), .C2(
        u1_srl_151_n144), .ZN(u1_srl_151_n138) );
  OAI211_X1 u1_srl_151_U146 ( .C1(u1_srl_151_n136), .C2(u1_srl_151_n96), .A(
        u1_srl_151_n137), .B(u1_srl_151_n138), .ZN(u1_adj_op_out_sft_9_) );
  INV_X4 u1_srl_151_U145 ( .A(u1_adj_op_10_), .ZN(u1_srl_151_n135) );
  INV_X4 u1_srl_151_U144 ( .A(u1_adj_op_11_), .ZN(u1_srl_151_n134) );
  INV_X4 u1_srl_151_U143 ( .A(n6261), .ZN(u1_srl_151_n133) );
  INV_X4 u1_srl_151_U142 ( .A(n6260), .ZN(u1_srl_151_n132) );
  INV_X4 u1_srl_151_U141 ( .A(n6259), .ZN(u1_srl_151_n131) );
  INV_X4 u1_srl_151_U140 ( .A(u1_adj_op_15_), .ZN(u1_srl_151_n130) );
  INV_X4 u1_srl_151_U139 ( .A(u1_adj_op_16_), .ZN(u1_srl_151_n129) );
  INV_X4 u1_srl_151_U138 ( .A(u1_adj_op_17_), .ZN(u1_srl_151_n128) );
  INV_X4 u1_srl_151_U137 ( .A(n6258), .ZN(u1_srl_151_n127) );
  INV_X4 u1_srl_151_U136 ( .A(n6257), .ZN(u1_srl_151_n126) );
  INV_X4 u1_srl_151_U135 ( .A(n6256), .ZN(u1_srl_151_n125) );
  INV_X4 u1_srl_151_U134 ( .A(u1_adj_op_20_), .ZN(u1_srl_151_n124) );
  INV_X4 u1_srl_151_U133 ( .A(u1_adj_op_21_), .ZN(u1_srl_151_n123) );
  INV_X4 u1_srl_151_U132 ( .A(u1_adj_op_22_), .ZN(u1_srl_151_n122) );
  INV_X4 u1_srl_151_U131 ( .A(n6255), .ZN(u1_srl_151_n121) );
  INV_X4 u1_srl_151_U130 ( .A(n6254), .ZN(u1_srl_151_n120) );
  INV_X4 u1_srl_151_U129 ( .A(n6253), .ZN(u1_srl_151_n119) );
  INV_X4 u1_srl_151_U128 ( .A(n6252), .ZN(u1_srl_151_n118) );
  INV_X4 u1_srl_151_U127 ( .A(u1_adj_op_27_), .ZN(u1_srl_151_n117) );
  INV_X4 u1_srl_151_U126 ( .A(u1_adj_op_28_), .ZN(u1_srl_151_n116) );
  INV_X4 u1_srl_151_U125 ( .A(n6251), .ZN(u1_srl_151_n115) );
  INV_X4 u1_srl_151_U124 ( .A(n6250), .ZN(u1_srl_151_n114) );
  INV_X4 u1_srl_151_U123 ( .A(n6249), .ZN(u1_srl_151_n113) );
  INV_X4 u1_srl_151_U122 ( .A(n6248), .ZN(u1_srl_151_n112) );
  INV_X4 u1_srl_151_U121 ( .A(u1_adj_op_32_), .ZN(u1_srl_151_n111) );
  INV_X4 u1_srl_151_U120 ( .A(n6247), .ZN(u1_srl_151_n110) );
  INV_X4 u1_srl_151_U119 ( .A(n6246), .ZN(u1_srl_151_n109) );
  INV_X4 u1_srl_151_U118 ( .A(n6245), .ZN(u1_srl_151_n108) );
  INV_X4 u1_srl_151_U117 ( .A(u1_adj_op_36_), .ZN(u1_srl_151_n107) );
  INV_X4 u1_srl_151_U116 ( .A(u1_adj_op_37_), .ZN(u1_srl_151_n106) );
  INV_X4 u1_srl_151_U115 ( .A(u1_adj_op_3_), .ZN(u1_srl_151_n105) );
  INV_X4 u1_srl_151_U114 ( .A(n6235), .ZN(u1_srl_151_n104) );
  INV_X4 u1_srl_151_U113 ( .A(n6233), .ZN(u1_srl_151_n103) );
  INV_X4 u1_srl_151_U112 ( .A(n6232), .ZN(u1_srl_151_n102) );
  INV_X4 u1_srl_151_U111 ( .A(n6231), .ZN(u1_srl_151_n101) );
  INV_X4 u1_srl_151_U110 ( .A(n6230), .ZN(u1_srl_151_n100) );
  INV_X4 u1_srl_151_U109 ( .A(n6229), .ZN(u1_srl_151_n99) );
  INV_X4 u1_srl_151_U108 ( .A(n6226), .ZN(u1_srl_151_n98) );
  INV_X4 u1_srl_151_U107 ( .A(n6225), .ZN(u1_srl_151_n97) );
  INV_X4 u1_srl_151_U106 ( .A(u1_srl_151_n145), .ZN(u1_srl_151_n95) );
  INV_X4 u1_srl_151_U105 ( .A(n6224), .ZN(u1_srl_151_n94) );
  INV_X4 u1_srl_151_U104 ( .A(n6222), .ZN(u1_srl_151_n93) );
  INV_X4 u1_srl_151_U103 ( .A(u1_srl_151_n302), .ZN(u1_srl_151_n92) );
  INV_X4 u1_srl_151_U102 ( .A(u1_srl_151_n266), .ZN(u1_srl_151_n91) );
  INV_X4 u1_srl_151_U101 ( .A(u1_srl_151_n178), .ZN(u1_srl_151_n90) );
  INV_X4 u1_srl_151_U100 ( .A(u1_srl_151_n303), .ZN(u1_srl_151_n89) );
  INV_X4 u1_srl_151_U99 ( .A(u1_srl_151_n233), .ZN(u1_srl_151_n88) );
  INV_X4 u1_srl_151_U98 ( .A(u1_srl_151_n238), .ZN(u1_srl_151_n87) );
  INV_X4 u1_srl_151_U97 ( .A(u1_srl_151_n306), .ZN(u1_srl_151_n86) );
  INV_X4 u1_srl_151_U96 ( .A(u1_srl_151_n267), .ZN(u1_srl_151_n85) );
  INV_X4 u1_srl_151_U95 ( .A(u1_srl_151_n161), .ZN(u1_srl_151_n84) );
  INV_X4 u1_srl_151_U94 ( .A(u1_srl_151_n319), .ZN(u1_srl_151_n83) );
  INV_X4 u1_srl_151_U93 ( .A(u1_srl_151_n320), .ZN(u1_srl_151_n82) );
  INV_X4 u1_srl_151_U92 ( .A(u1_srl_151_n321), .ZN(u1_srl_151_n81) );
  INV_X4 u1_srl_151_U91 ( .A(u1_srl_151_n254), .ZN(u1_srl_151_n80) );
  INV_X4 u1_srl_151_U90 ( .A(u1_srl_151_n281), .ZN(u1_srl_151_n79) );
  INV_X4 u1_srl_151_U89 ( .A(u1_srl_151_n324), .ZN(u1_srl_151_n78) );
  INV_X4 u1_srl_151_U88 ( .A(u1_srl_151_n283), .ZN(u1_srl_151_n77) );
  INV_X4 u1_srl_151_U87 ( .A(u1_srl_151_n248), .ZN(u1_srl_151_n76) );
  INV_X4 u1_srl_151_U86 ( .A(u1_srl_151_n279), .ZN(u1_srl_151_n75) );
  INV_X4 u1_srl_151_U85 ( .A(u1_srl_151_n334), .ZN(u1_srl_151_n74) );
  INV_X4 u1_srl_151_U84 ( .A(u1_srl_151_n262), .ZN(u1_srl_151_n73) );
  INV_X4 u1_srl_151_U83 ( .A(u1_srl_151_n177), .ZN(u1_srl_151_n72) );
  INV_X4 u1_srl_151_U82 ( .A(u1_srl_151_n335), .ZN(u1_srl_151_n71) );
  INV_X4 u1_srl_151_U81 ( .A(u1_srl_151_n286), .ZN(u1_srl_151_n70) );
  INV_X4 u1_srl_151_U80 ( .A(u1_srl_151_n336), .ZN(u1_srl_151_n69) );
  INV_X4 u1_srl_151_U79 ( .A(u1_srl_151_n263), .ZN(u1_srl_151_n68) );
  INV_X4 u1_srl_151_U78 ( .A(u1_srl_151_n348), .ZN(u1_srl_151_n67) );
  INV_X4 u1_srl_151_U77 ( .A(u1_srl_151_n179), .ZN(u1_srl_151_n66) );
  INV_X4 u1_srl_151_U76 ( .A(u1_srl_151_n349), .ZN(u1_srl_151_n65) );
  INV_X4 u1_srl_151_U75 ( .A(u1_srl_151_n241), .ZN(u1_srl_151_n64) );
  INV_X4 u1_srl_151_U74 ( .A(u1_srl_151_n351), .ZN(u1_srl_151_n63) );
  INV_X4 u1_srl_151_U73 ( .A(u1_srl_151_n312), .ZN(u1_srl_151_n62) );
  INV_X4 u1_srl_151_U72 ( .A(u1_srl_151_n352), .ZN(u1_srl_151_n61) );
  INV_X4 u1_srl_151_U71 ( .A(u1_srl_151_n270), .ZN(u1_srl_151_n60) );
  INV_X4 u1_srl_151_U70 ( .A(n6217), .ZN(u1_srl_151_n59) );
  INV_X4 u1_srl_151_U69 ( .A(u1_srl_151_n236), .ZN(u1_srl_151_n57) );
  INV_X4 u1_srl_151_U68 ( .A(u1_srl_151_n244), .ZN(u1_srl_151_n56) );
  INV_X4 u1_srl_151_U67 ( .A(u1_srl_151_n257), .ZN(u1_srl_151_n55) );
  INV_X4 u1_srl_151_U66 ( .A(u1_srl_151_n264), .ZN(u1_srl_151_n54) );
  INV_X4 u1_srl_151_U65 ( .A(u1_srl_151_n268), .ZN(u1_srl_151_n53) );
  INV_X4 u1_srl_151_U64 ( .A(u1_srl_151_n284), .ZN(u1_srl_151_n52) );
  INV_X4 u1_srl_151_U63 ( .A(u1_srl_151_n287), .ZN(u1_srl_151_n51) );
  INV_X4 u1_srl_151_U62 ( .A(u1_srl_151_n295), .ZN(u1_srl_151_n50) );
  INV_X4 u1_srl_151_U61 ( .A(u1_srl_151_n311), .ZN(u1_srl_151_n49) );
  INV_X4 u1_srl_151_U60 ( .A(u1_srl_151_n337), .ZN(u1_srl_151_n48) );
  INV_X4 u1_srl_151_U59 ( .A(u1_srl_151_n148), .ZN(u1_srl_151_n47) );
  INV_X4 u1_srl_151_U58 ( .A(u1_srl_151_n156), .ZN(u1_srl_151_n46) );
  INV_X4 u1_srl_151_U57 ( .A(u1_srl_151_n164), .ZN(u1_srl_151_n45) );
  INV_X4 u1_srl_151_U56 ( .A(u1_srl_151_n203), .ZN(u1_srl_151_n44) );
  INV_X4 u1_srl_151_U55 ( .A(u1_srl_151_n171), .ZN(u1_srl_151_n43) );
  INV_X4 u1_srl_151_U54 ( .A(u1_srl_151_n206), .ZN(u1_srl_151_n42) );
  INV_X4 u1_srl_151_U53 ( .A(u1_srl_151_n175), .ZN(u1_srl_151_n41) );
  INV_X4 u1_srl_151_U52 ( .A(u1_srl_151_n208), .ZN(u1_srl_151_n40) );
  INV_X4 u1_srl_151_U51 ( .A(u1_srl_151_n185), .ZN(u1_srl_151_n39) );
  INV_X4 u1_srl_151_U50 ( .A(u1_srl_151_n210), .ZN(u1_srl_151_n38) );
  INV_X4 u1_srl_151_U49 ( .A(u1_srl_151_n201), .ZN(u1_srl_151_n37) );
  INV_X4 u1_srl_151_U48 ( .A(u1_srl_151_n202), .ZN(u1_srl_151_n36) );
  INV_X4 u1_srl_151_U47 ( .A(u1_srl_151_n226), .ZN(u1_srl_151_n35) );
  INV_X4 u1_srl_151_U46 ( .A(u1_srl_151_n213), .ZN(u1_srl_151_n34) );
  INV_X4 u1_srl_151_U45 ( .A(u1_srl_151_n277), .ZN(u1_srl_151_n33) );
  INV_X4 u1_srl_151_U44 ( .A(u1_srl_151_n214), .ZN(u1_srl_151_n32) );
  INV_X4 u1_srl_151_U43 ( .A(u1_srl_151_n188), .ZN(u1_srl_151_n31) );
  INV_X4 u1_srl_151_U42 ( .A(u1_srl_151_n189), .ZN(u1_srl_151_n30) );
  INV_X4 u1_srl_151_U41 ( .A(u1_srl_151_n190), .ZN(u1_srl_151_n29) );
  INV_X4 u1_srl_151_U40 ( .A(u1_srl_151_n191), .ZN(u1_srl_151_n28) );
  INV_X4 u1_srl_151_U39 ( .A(u1_srl_151_n217), .ZN(u1_srl_151_n27) );
  INV_X4 u1_srl_151_U38 ( .A(u1_srl_151_n230), .ZN(u1_srl_151_n26) );
  INV_X4 u1_srl_151_U37 ( .A(u1_srl_151_n146), .ZN(u1_srl_151_n25) );
  INV_X4 u1_srl_151_U36 ( .A(u1_srl_151_n272), .ZN(u1_srl_151_n24) );
  INV_X4 u1_srl_151_U35 ( .A(u1_srl_151_n343), .ZN(u1_srl_151_n23) );
  INV_X4 u1_srl_151_U34 ( .A(u1_srl_151_n215), .ZN(u1_srl_151_n22) );
  INV_X4 u1_srl_151_U33 ( .A(u1_srl_151_n356), .ZN(u1_srl_151_n21) );
  INV_X4 u1_srl_151_U32 ( .A(u1_srl_151_n289), .ZN(u1_srl_151_n20) );
  INV_X4 u1_srl_151_U31 ( .A(u1_srl_151_n4), .ZN(u1_srl_151_n9) );
  INV_X4 u1_srl_151_U30 ( .A(u1_srl_151_n224), .ZN(u1_srl_151_n6) );
  INV_X4 u1_srl_151_U29 ( .A(u1_srl_151_n14), .ZN(u1_srl_151_n15) );
  INV_X4 u1_srl_151_U28 ( .A(u1_srl_151_n13), .ZN(u1_srl_151_n12) );
  INV_X4 u1_srl_151_U27 ( .A(u1_srl_151_n17), .ZN(u1_srl_151_n16) );
  INV_X4 u1_srl_151_U26 ( .A(u1_srl_151_n196), .ZN(u1_srl_151_n5) );
  NOR2_X2 u1_srl_151_U25 ( .A1(u1_srl_151_n1), .A2(u1_srl_151_n9), .ZN(
        u1_srl_151_n139) );
  INV_X4 u1_srl_151_U24 ( .A(u1_srl_151_n163), .ZN(u1_srl_151_n96) );
  INV_X4 u1_srl_151_U23 ( .A(u1_srl_151_n224), .ZN(u1_srl_151_n7) );
  INV_X4 u1_srl_151_U22 ( .A(u1_srl_151_n1), .ZN(u1_srl_151_n11) );
  INV_X4 u1_srl_151_U21 ( .A(u1_srl_151_n1), .ZN(u1_srl_151_n10) );
  INV_X4 u1_srl_151_U20 ( .A(u1_srl_151_n199), .ZN(u1_srl_151_n17) );
  INV_X4 u1_srl_151_U19 ( .A(u1_srl_151_n4), .ZN(u1_srl_151_n8) );
  INV_X4 u1_srl_151_U18 ( .A(u1_srl_151_n2), .ZN(u1_srl_151_n19) );
  NOR2_X2 u1_srl_151_U17 ( .A1(u1_srl_151_n94), .A2(n6217), .ZN(
        u1_srl_151_n196) );
  INV_X4 u1_srl_151_U16 ( .A(u1_srl_151_n198), .ZN(u1_srl_151_n14) );
  INV_X4 u1_srl_151_U15 ( .A(u1_srl_151_n3), .ZN(u1_srl_151_n13) );
  INV_X4 u1_srl_151_U14 ( .A(u1_srl_151_n19), .ZN(u1_srl_151_n18) );
  NOR2_X2 u1_srl_151_U13 ( .A1(u1_srl_151_n93), .A2(n6221), .ZN(
        u1_srl_151_n224) );
  AND2_X4 u1_srl_151_U12 ( .A1(u1_srl_151_n97), .A2(u1_srl_151_n98), .ZN(
        u1_srl_151_n4) );
  NAND2_X2 u1_srl_151_U11 ( .A1(n6221), .A2(u1_srl_151_n93), .ZN(u1_srl_151_n3) );
  NOR2_X2 u1_srl_151_U10 ( .A1(n6217), .A2(n6224), .ZN(u1_srl_151_n2) );
  OR2_X4 u1_srl_151_U9 ( .A1(u1_srl_151_n59), .A2(n6224), .ZN(u1_srl_151_n1)
         );
  NOR2_X2 u1_srl_151_U8 ( .A1(u1_srl_151_n98), .A2(n6225), .ZN(u1_srl_151_n145) );
  NOR2_X2 u1_srl_151_U7 ( .A1(u1_srl_151_n8), .A2(u1_srl_151_n58), .ZN(
        u1_srl_151_n141) );
  NOR2_X2 u1_srl_151_U6 ( .A1(u1_srl_151_n5), .A2(u1_srl_151_n8), .ZN(
        u1_srl_151_n143) );
  INV_X4 u1_srl_151_U5 ( .A(u1_srl_151_n237), .ZN(u1_srl_151_n58) );
  NOR2_X2 u1_srl_151_U4 ( .A1(u1_srl_151_n19), .A2(u1_srl_151_n8), .ZN(
        u1_srl_151_n146) );
  NOR2_X2 u1_srl_151_U3 ( .A1(u1_srl_151_n94), .A2(u1_srl_151_n59), .ZN(
        u1_srl_151_n237) );
  INV_X4 sub_1_root_u1_sub_133_aco_U12 ( .A(u1_N46), .ZN(
        sub_1_root_u1_sub_133_aco_n12) );
  INV_X4 sub_1_root_u1_sub_133_aco_U11 ( .A(u1_exp_small[0]), .ZN(
        sub_1_root_u1_sub_133_aco_n11) );
  INV_X4 sub_1_root_u1_sub_133_aco_U10 ( .A(u1_exp_small[10]), .ZN(
        sub_1_root_u1_sub_133_aco_n10) );
  INV_X4 sub_1_root_u1_sub_133_aco_U9 ( .A(u1_exp_small[1]), .ZN(
        sub_1_root_u1_sub_133_aco_n9) );
  INV_X4 sub_1_root_u1_sub_133_aco_U8 ( .A(u1_exp_small[2]), .ZN(
        sub_1_root_u1_sub_133_aco_n8) );
  INV_X4 sub_1_root_u1_sub_133_aco_U7 ( .A(u1_exp_small[3]), .ZN(
        sub_1_root_u1_sub_133_aco_n7) );
  INV_X4 sub_1_root_u1_sub_133_aco_U6 ( .A(u1_exp_small[4]), .ZN(
        sub_1_root_u1_sub_133_aco_n6) );
  INV_X4 sub_1_root_u1_sub_133_aco_U5 ( .A(u1_exp_small[5]), .ZN(
        sub_1_root_u1_sub_133_aco_n5) );
  INV_X4 sub_1_root_u1_sub_133_aco_U4 ( .A(u1_exp_small[6]), .ZN(
        sub_1_root_u1_sub_133_aco_n4) );
  INV_X4 sub_1_root_u1_sub_133_aco_U3 ( .A(u1_exp_small[7]), .ZN(
        sub_1_root_u1_sub_133_aco_n3) );
  INV_X4 sub_1_root_u1_sub_133_aco_U2 ( .A(n6228), .ZN(
        sub_1_root_u1_sub_133_aco_n2) );
  INV_X4 sub_1_root_u1_sub_133_aco_U1 ( .A(n6227), .ZN(
        sub_1_root_u1_sub_133_aco_n1) );
  FA_X1 sub_1_root_u1_sub_133_aco_U2_0 ( .A(u1_exp_large_0_), .B(
        sub_1_root_u1_sub_133_aco_n11), .CI(sub_1_root_u1_sub_133_aco_n12), 
        .CO(sub_1_root_u1_sub_133_aco_carry[1]), .S(u1_exp_diff2[0]) );
  FA_X1 sub_1_root_u1_sub_133_aco_U2_1 ( .A(u1_exp_large_1_), .B(
        sub_1_root_u1_sub_133_aco_n9), .CI(sub_1_root_u1_sub_133_aco_carry[1]), 
        .CO(sub_1_root_u1_sub_133_aco_carry[2]), .S(u1_exp_diff2[1]) );
  FA_X1 sub_1_root_u1_sub_133_aco_U2_2 ( .A(u1_exp_large_2_), .B(
        sub_1_root_u1_sub_133_aco_n8), .CI(sub_1_root_u1_sub_133_aco_carry[2]), 
        .CO(sub_1_root_u1_sub_133_aco_carry[3]), .S(u1_exp_diff2[2]) );
  FA_X1 sub_1_root_u1_sub_133_aco_U2_3 ( .A(u1_exp_large_3_), .B(
        sub_1_root_u1_sub_133_aco_n7), .CI(sub_1_root_u1_sub_133_aco_carry[3]), 
        .CO(sub_1_root_u1_sub_133_aco_carry[4]), .S(u1_exp_diff2[3]) );
  FA_X1 sub_1_root_u1_sub_133_aco_U2_4 ( .A(u1_exp_large_4_), .B(
        sub_1_root_u1_sub_133_aco_n6), .CI(sub_1_root_u1_sub_133_aco_carry[4]), 
        .CO(sub_1_root_u1_sub_133_aco_carry[5]), .S(u1_exp_diff2[4]) );
  FA_X1 sub_1_root_u1_sub_133_aco_U2_5 ( .A(u1_exp_large_5_), .B(
        sub_1_root_u1_sub_133_aco_n5), .CI(sub_1_root_u1_sub_133_aco_carry[5]), 
        .CO(sub_1_root_u1_sub_133_aco_carry[6]), .S(u1_exp_diff2[5]) );
  FA_X1 sub_1_root_u1_sub_133_aco_U2_6 ( .A(u1_exp_large_6_), .B(
        sub_1_root_u1_sub_133_aco_n4), .CI(sub_1_root_u1_sub_133_aco_carry[6]), 
        .CO(sub_1_root_u1_sub_133_aco_carry[7]), .S(u1_exp_diff2[6]) );
  FA_X1 sub_1_root_u1_sub_133_aco_U2_7 ( .A(u1_exp_large_7_), .B(
        sub_1_root_u1_sub_133_aco_n3), .CI(sub_1_root_u1_sub_133_aco_carry[7]), 
        .CO(sub_1_root_u1_sub_133_aco_carry[8]), .S(u1_exp_diff2[7]) );
  FA_X1 sub_1_root_u1_sub_133_aco_U2_8 ( .A(n6264), .B(
        sub_1_root_u1_sub_133_aco_n2), .CI(sub_1_root_u1_sub_133_aco_carry[8]), 
        .CO(sub_1_root_u1_sub_133_aco_carry[9]), .S(u1_exp_diff2[8]) );
  FA_X1 sub_1_root_u1_sub_133_aco_U2_9 ( .A(n6263), .B(
        sub_1_root_u1_sub_133_aco_n1), .CI(sub_1_root_u1_sub_133_aco_carry[9]), 
        .CO(sub_1_root_u1_sub_133_aco_carry[10]), .S(u1_exp_diff2[9]) );
  FA_X1 sub_1_root_u1_sub_133_aco_U2_10 ( .A(u1_exp_large_10_), .B(
        sub_1_root_u1_sub_133_aco_n10), .CI(
        sub_1_root_u1_sub_133_aco_carry[10]), .S(u1_exp_diff2[10]) );
  INV_X4 sub_436_3_U171 ( .A(N343), .ZN(sub_436_3_n171) );
  INV_X4 sub_436_3_U170 ( .A(opa_r1[1]), .ZN(sub_436_3_n170) );
  INV_X4 sub_436_3_U169 ( .A(opa_r1[2]), .ZN(sub_436_3_n169) );
  INV_X4 sub_436_3_U168 ( .A(opa_r1[3]), .ZN(sub_436_3_n168) );
  INV_X4 sub_436_3_U167 ( .A(opa_r1[4]), .ZN(sub_436_3_n167) );
  INV_X4 sub_436_3_U166 ( .A(opa_r1[5]), .ZN(sub_436_3_n166) );
  INV_X4 sub_436_3_U165 ( .A(opa_r1[6]), .ZN(sub_436_3_n165) );
  INV_X4 sub_436_3_U164 ( .A(opa_r1[7]), .ZN(sub_436_3_n164) );
  INV_X4 sub_436_3_U163 ( .A(opa_r1[8]), .ZN(sub_436_3_n163) );
  INV_X4 sub_436_3_U162 ( .A(opa_r1[9]), .ZN(sub_436_3_n162) );
  INV_X4 sub_436_3_U161 ( .A(opa_r1[10]), .ZN(sub_436_3_n161) );
  INV_X4 sub_436_3_U160 ( .A(opa_r1[11]), .ZN(sub_436_3_n160) );
  INV_X4 sub_436_3_U159 ( .A(opa_r1[12]), .ZN(sub_436_3_n159) );
  INV_X4 sub_436_3_U158 ( .A(opa_r1[13]), .ZN(sub_436_3_n158) );
  INV_X4 sub_436_3_U157 ( .A(opa_r1[14]), .ZN(sub_436_3_n157) );
  INV_X4 sub_436_3_U156 ( .A(opa_r1[15]), .ZN(sub_436_3_n156) );
  INV_X4 sub_436_3_U155 ( .A(opa_r1[16]), .ZN(sub_436_3_n155) );
  INV_X4 sub_436_3_U154 ( .A(opa_r1[17]), .ZN(sub_436_3_n154) );
  INV_X4 sub_436_3_U153 ( .A(opa_r1[18]), .ZN(sub_436_3_n153) );
  INV_X4 sub_436_3_U152 ( .A(opa_r1[19]), .ZN(sub_436_3_n152) );
  INV_X4 sub_436_3_U151 ( .A(opa_r1[20]), .ZN(sub_436_3_n151) );
  INV_X4 sub_436_3_U150 ( .A(opa_r1[21]), .ZN(sub_436_3_n150) );
  INV_X4 sub_436_3_U149 ( .A(opa_r1[22]), .ZN(sub_436_3_n149) );
  INV_X4 sub_436_3_U148 ( .A(opa_r1[23]), .ZN(sub_436_3_n148) );
  INV_X4 sub_436_3_U147 ( .A(opa_r1[24]), .ZN(sub_436_3_n147) );
  INV_X4 sub_436_3_U146 ( .A(opa_r1[25]), .ZN(sub_436_3_n146) );
  INV_X4 sub_436_3_U145 ( .A(opa_r1[26]), .ZN(sub_436_3_n145) );
  INV_X4 sub_436_3_U144 ( .A(opa_r1[27]), .ZN(sub_436_3_n144) );
  INV_X4 sub_436_3_U143 ( .A(opa_r1[28]), .ZN(sub_436_3_n143) );
  INV_X4 sub_436_3_U142 ( .A(opa_r1[29]), .ZN(sub_436_3_n142) );
  INV_X4 sub_436_3_U141 ( .A(opa_r1[30]), .ZN(sub_436_3_n141) );
  INV_X4 sub_436_3_U140 ( .A(opa_r1[31]), .ZN(sub_436_3_n140) );
  INV_X4 sub_436_3_U139 ( .A(opa_r1[32]), .ZN(sub_436_3_n139) );
  INV_X4 sub_436_3_U138 ( .A(opa_r1[33]), .ZN(sub_436_3_n138) );
  INV_X4 sub_436_3_U137 ( .A(opa_r1[34]), .ZN(sub_436_3_n137) );
  INV_X4 sub_436_3_U136 ( .A(opa_r1[35]), .ZN(sub_436_3_n136) );
  INV_X4 sub_436_3_U135 ( .A(opa_r1[36]), .ZN(sub_436_3_n135) );
  INV_X4 sub_436_3_U134 ( .A(opa_r1[37]), .ZN(sub_436_3_n134) );
  INV_X4 sub_436_3_U133 ( .A(opa_r1[38]), .ZN(sub_436_3_n133) );
  INV_X4 sub_436_3_U132 ( .A(opa_r1[39]), .ZN(sub_436_3_n132) );
  INV_X4 sub_436_3_U131 ( .A(opa_r1[40]), .ZN(sub_436_3_n131) );
  INV_X4 sub_436_3_U130 ( .A(opa_r1[41]), .ZN(sub_436_3_n130) );
  INV_X4 sub_436_3_U129 ( .A(opa_r1[42]), .ZN(sub_436_3_n129) );
  INV_X4 sub_436_3_U128 ( .A(opa_r1[43]), .ZN(sub_436_3_n128) );
  INV_X4 sub_436_3_U127 ( .A(opa_r1[44]), .ZN(sub_436_3_n127) );
  INV_X4 sub_436_3_U126 ( .A(opa_r1[45]), .ZN(sub_436_3_n126) );
  INV_X4 sub_436_3_U125 ( .A(opa_r1[46]), .ZN(sub_436_3_n125) );
  INV_X4 sub_436_3_U124 ( .A(opa_r1[47]), .ZN(sub_436_3_n124) );
  INV_X4 sub_436_3_U123 ( .A(opa_r1[48]), .ZN(sub_436_3_n123) );
  INV_X4 sub_436_3_U122 ( .A(opa_r1[49]), .ZN(sub_436_3_n122) );
  INV_X4 sub_436_3_U121 ( .A(opa_r1[50]), .ZN(sub_436_3_n121) );
  INV_X4 sub_436_3_U120 ( .A(opa_r1[51]), .ZN(sub_436_3_n120) );
  INV_X4 sub_436_3_U119 ( .A(opa_r1[52]), .ZN(sub_436_3_n119) );
  INV_X4 sub_436_3_U118 ( .A(opa_r1[53]), .ZN(sub_436_3_n118) );
  INV_X4 sub_436_3_U117 ( .A(opa_r1[54]), .ZN(sub_436_3_n117) );
  INV_X4 sub_436_3_U116 ( .A(opa_r1[55]), .ZN(sub_436_3_n116) );
  INV_X4 sub_436_3_U115 ( .A(opa_r1[56]), .ZN(sub_436_3_n115) );
  INV_X4 sub_436_3_U114 ( .A(opa_r1[57]), .ZN(sub_436_3_n114) );
  XOR2_X2 sub_436_3_U113 ( .A(sub_436_3_n158), .B(sub_436_3_n44), .Z(N513) );
  XOR2_X2 sub_436_3_U112 ( .A(sub_436_3_n159), .B(sub_436_3_n36), .Z(N512) );
  XOR2_X2 sub_436_3_U111 ( .A(sub_436_3_n160), .B(sub_436_3_n21), .Z(N511) );
  XOR2_X2 sub_436_3_U110 ( .A(sub_436_3_n161), .B(sub_436_3_n37), .Z(N510) );
  XOR2_X2 sub_436_3_U109 ( .A(sub_436_3_n162), .B(sub_436_3_n22), .Z(N509) );
  XOR2_X2 sub_436_3_U108 ( .A(sub_436_3_n164), .B(sub_436_3_n6), .Z(N507) );
  XOR2_X2 sub_436_3_U107 ( .A(sub_436_3_n168), .B(sub_436_3_n8), .Z(N503) );
  XOR2_X2 sub_436_3_U106 ( .A(sub_436_3_n169), .B(sub_436_3_n41), .Z(N502) );
  XOR2_X2 sub_436_3_U105 ( .A(sub_436_3_n163), .B(sub_436_3_n38), .Z(N508) );
  XOR2_X2 sub_436_3_U104 ( .A(sub_436_3_n165), .B(sub_436_3_n39), .Z(N506) );
  XOR2_X2 sub_436_3_U103 ( .A(sub_436_3_n166), .B(sub_436_3_n7), .Z(N505) );
  XOR2_X2 sub_436_3_U102 ( .A(sub_436_3_n167), .B(sub_436_3_n40), .Z(N504) );
  XOR2_X2 sub_436_3_U101 ( .A(sub_436_3_n170), .B(sub_436_3_n171), .Z(N501) );
  XOR2_X2 sub_436_3_U100 ( .A(sub_436_3_n117), .B(sub_436_3_n45), .Z(N554) );
  XOR2_X2 sub_436_3_U99 ( .A(sub_436_3_n118), .B(sub_436_3_n43), .Z(N553) );
  XOR2_X2 sub_436_3_U98 ( .A(sub_436_3_n119), .B(sub_436_3_n9), .Z(N552) );
  AND2_X4 sub_436_3_U97 ( .A1(sub_436_3_n115), .A2(sub_436_3_n46), .ZN(
        sub_436_3_n97) );
  XOR2_X2 sub_436_3_U96 ( .A(sub_436_3_n120), .B(sub_436_3_n42), .Z(N551) );
  AND2_X4 sub_436_3_U95 ( .A1(sub_436_3_n117), .A2(sub_436_3_n45), .ZN(
        sub_436_3_n95) );
  AND2_X4 sub_436_3_U94 ( .A1(sub_436_3_n158), .A2(sub_436_3_n44), .ZN(
        sub_436_3_n94) );
  AND2_X4 sub_436_3_U93 ( .A1(sub_436_3_n156), .A2(sub_436_3_n20), .ZN(
        sub_436_3_n93) );
  AND2_X4 sub_436_3_U92 ( .A1(sub_436_3_n154), .A2(sub_436_3_n19), .ZN(
        sub_436_3_n92) );
  AND2_X4 sub_436_3_U91 ( .A1(sub_436_3_n152), .A2(sub_436_3_n18), .ZN(
        sub_436_3_n91) );
  AND2_X4 sub_436_3_U90 ( .A1(sub_436_3_n150), .A2(sub_436_3_n17), .ZN(
        sub_436_3_n90) );
  AND2_X4 sub_436_3_U89 ( .A1(sub_436_3_n148), .A2(sub_436_3_n52), .ZN(
        sub_436_3_n89) );
  AND2_X4 sub_436_3_U88 ( .A1(sub_436_3_n146), .A2(sub_436_3_n51), .ZN(
        sub_436_3_n88) );
  AND2_X4 sub_436_3_U87 ( .A1(sub_436_3_n144), .A2(sub_436_3_n50), .ZN(
        sub_436_3_n87) );
  AND2_X4 sub_436_3_U86 ( .A1(sub_436_3_n142), .A2(sub_436_3_n49), .ZN(
        sub_436_3_n86) );
  AND2_X4 sub_436_3_U85 ( .A1(sub_436_3_n140), .A2(sub_436_3_n48), .ZN(
        sub_436_3_n85) );
  AND2_X4 sub_436_3_U84 ( .A1(sub_436_3_n138), .A2(sub_436_3_n23), .ZN(
        sub_436_3_n84) );
  AND2_X4 sub_436_3_U83 ( .A1(sub_436_3_n136), .A2(sub_436_3_n16), .ZN(
        sub_436_3_n83) );
  AND2_X4 sub_436_3_U82 ( .A1(sub_436_3_n134), .A2(sub_436_3_n15), .ZN(
        sub_436_3_n82) );
  AND2_X4 sub_436_3_U81 ( .A1(sub_436_3_n132), .A2(sub_436_3_n14), .ZN(
        sub_436_3_n81) );
  AND2_X4 sub_436_3_U80 ( .A1(sub_436_3_n130), .A2(sub_436_3_n13), .ZN(
        sub_436_3_n80) );
  AND2_X4 sub_436_3_U79 ( .A1(sub_436_3_n128), .A2(sub_436_3_n12), .ZN(
        sub_436_3_n79) );
  AND2_X4 sub_436_3_U78 ( .A1(sub_436_3_n126), .A2(sub_436_3_n11), .ZN(
        sub_436_3_n78) );
  AND2_X4 sub_436_3_U77 ( .A1(sub_436_3_n124), .A2(sub_436_3_n10), .ZN(
        sub_436_3_n77) );
  AND2_X4 sub_436_3_U76 ( .A1(sub_436_3_n122), .A2(sub_436_3_n47), .ZN(
        sub_436_3_n76) );
  XOR2_X2 sub_436_3_U75 ( .A(sub_436_3_n150), .B(sub_436_3_n17), .Z(N521) );
  XOR2_X2 sub_436_3_U74 ( .A(sub_436_3_n151), .B(sub_436_3_n91), .Z(N520) );
  XOR2_X2 sub_436_3_U73 ( .A(sub_436_3_n156), .B(sub_436_3_n20), .Z(N515) );
  XOR2_X2 sub_436_3_U72 ( .A(sub_436_3_n157), .B(sub_436_3_n94), .Z(N514) );
  XOR2_X2 sub_436_3_U71 ( .A(sub_436_3_n152), .B(sub_436_3_n18), .Z(N519) );
  XOR2_X2 sub_436_3_U70 ( .A(sub_436_3_n153), .B(sub_436_3_n92), .Z(N518) );
  XOR2_X2 sub_436_3_U69 ( .A(sub_436_3_n154), .B(sub_436_3_n19), .Z(N517) );
  XOR2_X2 sub_436_3_U68 ( .A(sub_436_3_n155), .B(sub_436_3_n93), .Z(N516) );
  XOR2_X2 sub_436_3_U67 ( .A(sub_436_3_n124), .B(sub_436_3_n10), .Z(N547) );
  XOR2_X2 sub_436_3_U66 ( .A(sub_436_3_n125), .B(sub_436_3_n78), .Z(N546) );
  XOR2_X2 sub_436_3_U65 ( .A(sub_436_3_n126), .B(sub_436_3_n11), .Z(N545) );
  XOR2_X2 sub_436_3_U64 ( .A(sub_436_3_n127), .B(sub_436_3_n79), .Z(N544) );
  XOR2_X2 sub_436_3_U63 ( .A(sub_436_3_n128), .B(sub_436_3_n12), .Z(N543) );
  XOR2_X2 sub_436_3_U62 ( .A(sub_436_3_n130), .B(sub_436_3_n13), .Z(N541) );
  XOR2_X2 sub_436_3_U61 ( .A(sub_436_3_n132), .B(sub_436_3_n14), .Z(N539) );
  XOR2_X2 sub_436_3_U60 ( .A(sub_436_3_n133), .B(sub_436_3_n82), .Z(N538) );
  XOR2_X2 sub_436_3_U59 ( .A(sub_436_3_n134), .B(sub_436_3_n15), .Z(N537) );
  XOR2_X2 sub_436_3_U58 ( .A(sub_436_3_n135), .B(sub_436_3_n83), .Z(N536) );
  XOR2_X2 sub_436_3_U57 ( .A(sub_436_3_n138), .B(sub_436_3_n23), .Z(N533) );
  XOR2_X2 sub_436_3_U56 ( .A(sub_436_3_n129), .B(sub_436_3_n80), .Z(N542) );
  XOR2_X2 sub_436_3_U55 ( .A(sub_436_3_n131), .B(sub_436_3_n81), .Z(N540) );
  XOR2_X2 sub_436_3_U54 ( .A(sub_436_3_n136), .B(sub_436_3_n16), .Z(N535) );
  XOR2_X2 sub_436_3_U53 ( .A(sub_436_3_n137), .B(sub_436_3_n84), .Z(N534) );
  AND2_X4 sub_436_3_U52 ( .A1(sub_436_3_n149), .A2(sub_436_3_n90), .ZN(
        sub_436_3_n52) );
  AND2_X4 sub_436_3_U51 ( .A1(sub_436_3_n147), .A2(sub_436_3_n89), .ZN(
        sub_436_3_n51) );
  AND2_X4 sub_436_3_U50 ( .A1(sub_436_3_n145), .A2(sub_436_3_n88), .ZN(
        sub_436_3_n50) );
  AND2_X4 sub_436_3_U49 ( .A1(sub_436_3_n143), .A2(sub_436_3_n87), .ZN(
        sub_436_3_n49) );
  AND2_X4 sub_436_3_U48 ( .A1(sub_436_3_n141), .A2(sub_436_3_n86), .ZN(
        sub_436_3_n48) );
  AND2_X4 sub_436_3_U47 ( .A1(sub_436_3_n123), .A2(sub_436_3_n77), .ZN(
        sub_436_3_n47) );
  AND2_X4 sub_436_3_U46 ( .A1(sub_436_3_n116), .A2(sub_436_3_n95), .ZN(
        sub_436_3_n46) );
  AND2_X4 sub_436_3_U45 ( .A1(sub_436_3_n118), .A2(sub_436_3_n43), .ZN(
        sub_436_3_n45) );
  AND2_X4 sub_436_3_U44 ( .A1(sub_436_3_n159), .A2(sub_436_3_n36), .ZN(
        sub_436_3_n44) );
  AND2_X4 sub_436_3_U43 ( .A1(sub_436_3_n119), .A2(sub_436_3_n9), .ZN(
        sub_436_3_n43) );
  AND2_X4 sub_436_3_U42 ( .A1(sub_436_3_n121), .A2(sub_436_3_n76), .ZN(
        sub_436_3_n42) );
  AND2_X4 sub_436_3_U41 ( .A1(sub_436_3_n170), .A2(sub_436_3_n171), .ZN(
        sub_436_3_n41) );
  AND2_X4 sub_436_3_U40 ( .A1(sub_436_3_n168), .A2(sub_436_3_n8), .ZN(
        sub_436_3_n40) );
  AND2_X4 sub_436_3_U39 ( .A1(sub_436_3_n166), .A2(sub_436_3_n7), .ZN(
        sub_436_3_n39) );
  AND2_X4 sub_436_3_U38 ( .A1(sub_436_3_n164), .A2(sub_436_3_n6), .ZN(
        sub_436_3_n38) );
  AND2_X4 sub_436_3_U37 ( .A1(sub_436_3_n162), .A2(sub_436_3_n22), .ZN(
        sub_436_3_n37) );
  AND2_X4 sub_436_3_U36 ( .A1(sub_436_3_n160), .A2(sub_436_3_n21), .ZN(
        sub_436_3_n36) );
  XOR2_X2 sub_436_3_U35 ( .A(sub_436_3_n144), .B(sub_436_3_n50), .Z(N527) );
  XOR2_X2 sub_436_3_U34 ( .A(sub_436_3_n145), .B(sub_436_3_n88), .Z(N526) );
  XOR2_X2 sub_436_3_U33 ( .A(sub_436_3_n146), .B(sub_436_3_n51), .Z(N525) );
  XOR2_X2 sub_436_3_U32 ( .A(sub_436_3_n148), .B(sub_436_3_n52), .Z(N523) );
  XOR2_X2 sub_436_3_U31 ( .A(sub_436_3_n149), .B(sub_436_3_n90), .Z(N522) );
  XOR2_X2 sub_436_3_U30 ( .A(sub_436_3_n143), .B(sub_436_3_n87), .Z(N528) );
  XOR2_X2 sub_436_3_U29 ( .A(sub_436_3_n147), .B(sub_436_3_n89), .Z(N524) );
  XOR2_X2 sub_436_3_U28 ( .A(sub_436_3_n141), .B(sub_436_3_n86), .Z(N530) );
  XOR2_X2 sub_436_3_U27 ( .A(sub_436_3_n142), .B(sub_436_3_n49), .Z(N529) );
  XOR2_X2 sub_436_3_U26 ( .A(sub_436_3_n121), .B(sub_436_3_n76), .Z(N550) );
  XOR2_X2 sub_436_3_U25 ( .A(sub_436_3_n123), .B(sub_436_3_n77), .Z(N548) );
  XOR2_X2 sub_436_3_U24 ( .A(sub_436_3_n122), .B(sub_436_3_n47), .Z(N549) );
  AND2_X4 sub_436_3_U23 ( .A1(sub_436_3_n139), .A2(sub_436_3_n85), .ZN(
        sub_436_3_n23) );
  AND2_X4 sub_436_3_U22 ( .A1(sub_436_3_n163), .A2(sub_436_3_n38), .ZN(
        sub_436_3_n22) );
  AND2_X4 sub_436_3_U21 ( .A1(sub_436_3_n161), .A2(sub_436_3_n37), .ZN(
        sub_436_3_n21) );
  AND2_X4 sub_436_3_U20 ( .A1(sub_436_3_n157), .A2(sub_436_3_n94), .ZN(
        sub_436_3_n20) );
  AND2_X4 sub_436_3_U19 ( .A1(sub_436_3_n155), .A2(sub_436_3_n93), .ZN(
        sub_436_3_n19) );
  AND2_X4 sub_436_3_U18 ( .A1(sub_436_3_n153), .A2(sub_436_3_n92), .ZN(
        sub_436_3_n18) );
  AND2_X4 sub_436_3_U17 ( .A1(sub_436_3_n151), .A2(sub_436_3_n91), .ZN(
        sub_436_3_n17) );
  AND2_X4 sub_436_3_U16 ( .A1(sub_436_3_n137), .A2(sub_436_3_n84), .ZN(
        sub_436_3_n16) );
  AND2_X4 sub_436_3_U15 ( .A1(sub_436_3_n135), .A2(sub_436_3_n83), .ZN(
        sub_436_3_n15) );
  AND2_X4 sub_436_3_U14 ( .A1(sub_436_3_n133), .A2(sub_436_3_n82), .ZN(
        sub_436_3_n14) );
  AND2_X4 sub_436_3_U13 ( .A1(sub_436_3_n131), .A2(sub_436_3_n81), .ZN(
        sub_436_3_n13) );
  AND2_X4 sub_436_3_U12 ( .A1(sub_436_3_n129), .A2(sub_436_3_n80), .ZN(
        sub_436_3_n12) );
  AND2_X4 sub_436_3_U11 ( .A1(sub_436_3_n127), .A2(sub_436_3_n79), .ZN(
        sub_436_3_n11) );
  AND2_X4 sub_436_3_U10 ( .A1(sub_436_3_n125), .A2(sub_436_3_n78), .ZN(
        sub_436_3_n10) );
  AND2_X4 sub_436_3_U9 ( .A1(sub_436_3_n120), .A2(sub_436_3_n42), .ZN(
        sub_436_3_n9) );
  AND2_X4 sub_436_3_U8 ( .A1(sub_436_3_n169), .A2(sub_436_3_n41), .ZN(
        sub_436_3_n8) );
  AND2_X4 sub_436_3_U7 ( .A1(sub_436_3_n167), .A2(sub_436_3_n40), .ZN(
        sub_436_3_n7) );
  AND2_X4 sub_436_3_U6 ( .A1(sub_436_3_n165), .A2(sub_436_3_n39), .ZN(
        sub_436_3_n6) );
  XOR2_X2 sub_436_3_U5 ( .A(sub_436_3_n139), .B(sub_436_3_n85), .Z(N532) );
  XOR2_X2 sub_436_3_U4 ( .A(sub_436_3_n140), .B(sub_436_3_n48), .Z(N531) );
  XOR2_X2 sub_436_3_U3 ( .A(sub_436_3_n114), .B(sub_436_3_n97), .Z(N557) );
  XOR2_X2 sub_436_3_U2 ( .A(sub_436_3_n115), .B(sub_436_3_n46), .Z(N556) );
  XOR2_X2 sub_436_3_U1 ( .A(sub_436_3_n116), .B(sub_436_3_n95), .Z(N555) );
  INV_X4 sub_436_b0_U157 ( .A(N343), .ZN(sub_436_b0_n157) );
  INV_X4 sub_436_b0_U156 ( .A(opa_r1[1]), .ZN(sub_436_b0_n156) );
  INV_X4 sub_436_b0_U155 ( .A(opa_r1[2]), .ZN(sub_436_b0_n155) );
  INV_X4 sub_436_b0_U154 ( .A(opa_r1[3]), .ZN(sub_436_b0_n154) );
  INV_X4 sub_436_b0_U153 ( .A(opa_r1[4]), .ZN(sub_436_b0_n153) );
  INV_X4 sub_436_b0_U152 ( .A(opa_r1[5]), .ZN(sub_436_b0_n152) );
  INV_X4 sub_436_b0_U151 ( .A(opa_r1[6]), .ZN(sub_436_b0_n151) );
  INV_X4 sub_436_b0_U150 ( .A(opa_r1[7]), .ZN(sub_436_b0_n150) );
  INV_X4 sub_436_b0_U149 ( .A(opa_r1[8]), .ZN(sub_436_b0_n149) );
  INV_X4 sub_436_b0_U148 ( .A(opa_r1[9]), .ZN(sub_436_b0_n148) );
  INV_X4 sub_436_b0_U147 ( .A(opa_r1[10]), .ZN(sub_436_b0_n147) );
  INV_X4 sub_436_b0_U146 ( .A(opa_r1[11]), .ZN(sub_436_b0_n146) );
  INV_X4 sub_436_b0_U145 ( .A(opa_r1[12]), .ZN(sub_436_b0_n145) );
  INV_X4 sub_436_b0_U144 ( .A(opa_r1[13]), .ZN(sub_436_b0_n144) );
  INV_X4 sub_436_b0_U143 ( .A(opa_r1[14]), .ZN(sub_436_b0_n143) );
  INV_X4 sub_436_b0_U142 ( .A(opa_r1[15]), .ZN(sub_436_b0_n142) );
  INV_X4 sub_436_b0_U141 ( .A(opa_r1[16]), .ZN(sub_436_b0_n141) );
  INV_X4 sub_436_b0_U140 ( .A(opa_r1[17]), .ZN(sub_436_b0_n140) );
  INV_X4 sub_436_b0_U139 ( .A(opa_r1[18]), .ZN(sub_436_b0_n139) );
  INV_X4 sub_436_b0_U138 ( .A(opa_r1[19]), .ZN(sub_436_b0_n138) );
  INV_X4 sub_436_b0_U137 ( .A(opa_r1[20]), .ZN(sub_436_b0_n137) );
  INV_X4 sub_436_b0_U136 ( .A(opa_r1[21]), .ZN(sub_436_b0_n136) );
  INV_X4 sub_436_b0_U135 ( .A(opa_r1[22]), .ZN(sub_436_b0_n135) );
  INV_X4 sub_436_b0_U134 ( .A(opa_r1[23]), .ZN(sub_436_b0_n134) );
  INV_X4 sub_436_b0_U133 ( .A(opa_r1[24]), .ZN(sub_436_b0_n133) );
  INV_X4 sub_436_b0_U132 ( .A(opa_r1[25]), .ZN(sub_436_b0_n132) );
  INV_X4 sub_436_b0_U131 ( .A(opa_r1[26]), .ZN(sub_436_b0_n131) );
  INV_X4 sub_436_b0_U130 ( .A(opa_r1[27]), .ZN(sub_436_b0_n130) );
  INV_X4 sub_436_b0_U129 ( .A(opa_r1[28]), .ZN(sub_436_b0_n129) );
  INV_X4 sub_436_b0_U128 ( .A(opa_r1[29]), .ZN(sub_436_b0_n128) );
  INV_X4 sub_436_b0_U127 ( .A(opa_r1[30]), .ZN(sub_436_b0_n127) );
  INV_X4 sub_436_b0_U126 ( .A(opa_r1[31]), .ZN(sub_436_b0_n126) );
  INV_X4 sub_436_b0_U125 ( .A(opa_r1[32]), .ZN(sub_436_b0_n125) );
  INV_X4 sub_436_b0_U124 ( .A(opa_r1[33]), .ZN(sub_436_b0_n124) );
  INV_X4 sub_436_b0_U123 ( .A(opa_r1[34]), .ZN(sub_436_b0_n123) );
  INV_X4 sub_436_b0_U122 ( .A(opa_r1[35]), .ZN(sub_436_b0_n122) );
  INV_X4 sub_436_b0_U121 ( .A(opa_r1[36]), .ZN(sub_436_b0_n121) );
  INV_X4 sub_436_b0_U120 ( .A(opa_r1[37]), .ZN(sub_436_b0_n120) );
  INV_X4 sub_436_b0_U119 ( .A(opa_r1[38]), .ZN(sub_436_b0_n119) );
  INV_X4 sub_436_b0_U118 ( .A(opa_r1[39]), .ZN(sub_436_b0_n118) );
  INV_X4 sub_436_b0_U117 ( .A(opa_r1[40]), .ZN(sub_436_b0_n117) );
  INV_X4 sub_436_b0_U116 ( .A(opa_r1[41]), .ZN(sub_436_b0_n116) );
  INV_X4 sub_436_b0_U115 ( .A(opa_r1[42]), .ZN(sub_436_b0_n115) );
  INV_X4 sub_436_b0_U114 ( .A(opa_r1[43]), .ZN(sub_436_b0_n114) );
  INV_X4 sub_436_b0_U113 ( .A(opa_r1[44]), .ZN(sub_436_b0_n113) );
  INV_X4 sub_436_b0_U112 ( .A(opa_r1[45]), .ZN(sub_436_b0_n112) );
  INV_X4 sub_436_b0_U111 ( .A(opa_r1[46]), .ZN(sub_436_b0_n111) );
  INV_X4 sub_436_b0_U110 ( .A(opa_r1[47]), .ZN(sub_436_b0_n110) );
  INV_X4 sub_436_b0_U109 ( .A(opa_r1[48]), .ZN(sub_436_b0_n109) );
  INV_X4 sub_436_b0_U108 ( .A(opa_r1[49]), .ZN(sub_436_b0_n108) );
  INV_X4 sub_436_b0_U107 ( .A(opa_r1[50]), .ZN(sub_436_b0_n107) );
  INV_X4 sub_436_b0_U106 ( .A(opa_r1[51]), .ZN(sub_436_b0_n106) );
  INV_X4 sub_436_b0_U105 ( .A(N340), .ZN(sub_436_b0_n105) );
  NAND2_X2 sub_436_b0_U104 ( .A1(sub_436_b0_n105), .A2(sub_436_b0_n1), .ZN(
        N396) );
  XOR2_X2 sub_436_b0_U103 ( .A(sub_436_b0_n144), .B(sub_436_b0_n12), .Z(N356)
         );
  XOR2_X2 sub_436_b0_U102 ( .A(sub_436_b0_n145), .B(sub_436_b0_n63), .Z(N355)
         );
  XOR2_X2 sub_436_b0_U101 ( .A(sub_436_b0_n146), .B(sub_436_b0_n13), .Z(N354)
         );
  XOR2_X2 sub_436_b0_U100 ( .A(sub_436_b0_n147), .B(sub_436_b0_n64), .Z(N353)
         );
  XOR2_X2 sub_436_b0_U99 ( .A(sub_436_b0_n148), .B(sub_436_b0_n14), .Z(N352)
         );
  XOR2_X2 sub_436_b0_U98 ( .A(sub_436_b0_n149), .B(sub_436_b0_n65), .Z(N351)
         );
  XOR2_X2 sub_436_b0_U97 ( .A(sub_436_b0_n150), .B(sub_436_b0_n15), .Z(N350)
         );
  XOR2_X2 sub_436_b0_U96 ( .A(sub_436_b0_n122), .B(sub_436_b0_n17), .Z(N378)
         );
  XOR2_X2 sub_436_b0_U95 ( .A(sub_436_b0_n123), .B(sub_436_b0_n52), .Z(N377)
         );
  XOR2_X2 sub_436_b0_U94 ( .A(sub_436_b0_n124), .B(sub_436_b0_n18), .Z(N376)
         );
  XOR2_X2 sub_436_b0_U93 ( .A(sub_436_b0_n125), .B(sub_436_b0_n53), .Z(N375)
         );
  XOR2_X2 sub_436_b0_U92 ( .A(sub_436_b0_n126), .B(sub_436_b0_n19), .Z(N374)
         );
  XOR2_X2 sub_436_b0_U91 ( .A(sub_436_b0_n127), .B(sub_436_b0_n54), .Z(N373)
         );
  XOR2_X2 sub_436_b0_U90 ( .A(sub_436_b0_n128), .B(sub_436_b0_n20), .Z(N372)
         );
  XOR2_X2 sub_436_b0_U89 ( .A(sub_436_b0_n129), .B(sub_436_b0_n55), .Z(N371)
         );
  XOR2_X2 sub_436_b0_U88 ( .A(sub_436_b0_n130), .B(sub_436_b0_n21), .Z(N370)
         );
  XOR2_X2 sub_436_b0_U87 ( .A(sub_436_b0_n131), .B(sub_436_b0_n56), .Z(N369)
         );
  XOR2_X2 sub_436_b0_U86 ( .A(sub_436_b0_n132), .B(sub_436_b0_n22), .Z(N368)
         );
  XOR2_X2 sub_436_b0_U85 ( .A(sub_436_b0_n133), .B(sub_436_b0_n57), .Z(N367)
         );
  XOR2_X2 sub_436_b0_U84 ( .A(sub_436_b0_n134), .B(sub_436_b0_n23), .Z(N366)
         );
  XOR2_X2 sub_436_b0_U83 ( .A(sub_436_b0_n135), .B(sub_436_b0_n58), .Z(N365)
         );
  XOR2_X2 sub_436_b0_U82 ( .A(sub_436_b0_n136), .B(sub_436_b0_n24), .Z(N364)
         );
  XOR2_X2 sub_436_b0_U81 ( .A(sub_436_b0_n137), .B(sub_436_b0_n59), .Z(N363)
         );
  XOR2_X2 sub_436_b0_U80 ( .A(sub_436_b0_n138), .B(sub_436_b0_n25), .Z(N362)
         );
  XOR2_X2 sub_436_b0_U79 ( .A(sub_436_b0_n139), .B(sub_436_b0_n60), .Z(N361)
         );
  XOR2_X2 sub_436_b0_U78 ( .A(sub_436_b0_n140), .B(sub_436_b0_n26), .Z(N360)
         );
  XOR2_X2 sub_436_b0_U77 ( .A(sub_436_b0_n141), .B(sub_436_b0_n61), .Z(N359)
         );
  XOR2_X2 sub_436_b0_U76 ( .A(sub_436_b0_n142), .B(sub_436_b0_n11), .Z(N358)
         );
  XOR2_X2 sub_436_b0_U75 ( .A(sub_436_b0_n143), .B(sub_436_b0_n62), .Z(N357)
         );
  XOR2_X2 sub_436_b0_U74 ( .A(sub_436_b0_n105), .B(sub_436_b0_n1), .Z(N395) );
  XOR2_X2 sub_436_b0_U73 ( .A(sub_436_b0_n106), .B(sub_436_b0_n10), .Z(N394)
         );
  XOR2_X2 sub_436_b0_U72 ( .A(sub_436_b0_n108), .B(sub_436_b0_n27), .Z(N392)
         );
  XOR2_X2 sub_436_b0_U71 ( .A(sub_436_b0_n110), .B(sub_436_b0_n16), .Z(N390)
         );
  XOR2_X2 sub_436_b0_U70 ( .A(sub_436_b0_n111), .B(sub_436_b0_n46), .Z(N389)
         );
  XOR2_X2 sub_436_b0_U69 ( .A(sub_436_b0_n121), .B(sub_436_b0_n51), .Z(N379)
         );
  AND2_X4 sub_436_b0_U68 ( .A1(sub_436_b0_n156), .A2(sub_436_b0_n157), .ZN(
        sub_436_b0_n68) );
  AND2_X4 sub_436_b0_U67 ( .A1(sub_436_b0_n154), .A2(sub_436_b0_n30), .ZN(
        sub_436_b0_n67) );
  AND2_X4 sub_436_b0_U66 ( .A1(sub_436_b0_n152), .A2(sub_436_b0_n28), .ZN(
        sub_436_b0_n66) );
  AND2_X4 sub_436_b0_U65 ( .A1(sub_436_b0_n150), .A2(sub_436_b0_n15), .ZN(
        sub_436_b0_n65) );
  AND2_X4 sub_436_b0_U64 ( .A1(sub_436_b0_n148), .A2(sub_436_b0_n14), .ZN(
        sub_436_b0_n64) );
  AND2_X4 sub_436_b0_U63 ( .A1(sub_436_b0_n146), .A2(sub_436_b0_n13), .ZN(
        sub_436_b0_n63) );
  AND2_X4 sub_436_b0_U62 ( .A1(sub_436_b0_n144), .A2(sub_436_b0_n12), .ZN(
        sub_436_b0_n62) );
  AND2_X4 sub_436_b0_U61 ( .A1(sub_436_b0_n142), .A2(sub_436_b0_n11), .ZN(
        sub_436_b0_n61) );
  AND2_X4 sub_436_b0_U60 ( .A1(sub_436_b0_n140), .A2(sub_436_b0_n26), .ZN(
        sub_436_b0_n60) );
  AND2_X4 sub_436_b0_U59 ( .A1(sub_436_b0_n138), .A2(sub_436_b0_n25), .ZN(
        sub_436_b0_n59) );
  AND2_X4 sub_436_b0_U58 ( .A1(sub_436_b0_n136), .A2(sub_436_b0_n24), .ZN(
        sub_436_b0_n58) );
  AND2_X4 sub_436_b0_U57 ( .A1(sub_436_b0_n134), .A2(sub_436_b0_n23), .ZN(
        sub_436_b0_n57) );
  AND2_X4 sub_436_b0_U56 ( .A1(sub_436_b0_n132), .A2(sub_436_b0_n22), .ZN(
        sub_436_b0_n56) );
  AND2_X4 sub_436_b0_U55 ( .A1(sub_436_b0_n130), .A2(sub_436_b0_n21), .ZN(
        sub_436_b0_n55) );
  AND2_X4 sub_436_b0_U54 ( .A1(sub_436_b0_n128), .A2(sub_436_b0_n20), .ZN(
        sub_436_b0_n54) );
  AND2_X4 sub_436_b0_U53 ( .A1(sub_436_b0_n126), .A2(sub_436_b0_n19), .ZN(
        sub_436_b0_n53) );
  AND2_X4 sub_436_b0_U52 ( .A1(sub_436_b0_n124), .A2(sub_436_b0_n18), .ZN(
        sub_436_b0_n52) );
  AND2_X4 sub_436_b0_U51 ( .A1(sub_436_b0_n122), .A2(sub_436_b0_n17), .ZN(
        sub_436_b0_n51) );
  AND2_X4 sub_436_b0_U50 ( .A1(sub_436_b0_n120), .A2(sub_436_b0_n29), .ZN(
        sub_436_b0_n50) );
  AND2_X4 sub_436_b0_U49 ( .A1(sub_436_b0_n118), .A2(sub_436_b0_n34), .ZN(
        sub_436_b0_n49) );
  AND2_X4 sub_436_b0_U48 ( .A1(sub_436_b0_n116), .A2(sub_436_b0_n33), .ZN(
        sub_436_b0_n48) );
  AND2_X4 sub_436_b0_U47 ( .A1(sub_436_b0_n114), .A2(sub_436_b0_n32), .ZN(
        sub_436_b0_n47) );
  AND2_X4 sub_436_b0_U46 ( .A1(sub_436_b0_n112), .A2(sub_436_b0_n31), .ZN(
        sub_436_b0_n46) );
  AND2_X4 sub_436_b0_U45 ( .A1(sub_436_b0_n110), .A2(sub_436_b0_n16), .ZN(
        sub_436_b0_n45) );
  AND2_X4 sub_436_b0_U44 ( .A1(sub_436_b0_n108), .A2(sub_436_b0_n27), .ZN(
        sub_436_b0_n44) );
  XOR2_X2 sub_436_b0_U43 ( .A(sub_436_b0_n151), .B(sub_436_b0_n66), .Z(N349)
         );
  XOR2_X2 sub_436_b0_U42 ( .A(sub_436_b0_n152), .B(sub_436_b0_n28), .Z(N348)
         );
  XOR2_X2 sub_436_b0_U41 ( .A(sub_436_b0_n153), .B(sub_436_b0_n67), .Z(N347)
         );
  XOR2_X2 sub_436_b0_U40 ( .A(sub_436_b0_n154), .B(sub_436_b0_n30), .Z(N346)
         );
  XOR2_X2 sub_436_b0_U39 ( .A(sub_436_b0_n155), .B(sub_436_b0_n68), .Z(N345)
         );
  XOR2_X2 sub_436_b0_U38 ( .A(sub_436_b0_n156), .B(sub_436_b0_n157), .Z(N344)
         );
  XOR2_X2 sub_436_b0_U37 ( .A(sub_436_b0_n109), .B(sub_436_b0_n45), .Z(N391)
         );
  XOR2_X2 sub_436_b0_U36 ( .A(sub_436_b0_n112), .B(sub_436_b0_n31), .Z(N388)
         );
  XOR2_X2 sub_436_b0_U35 ( .A(sub_436_b0_n107), .B(sub_436_b0_n44), .Z(N393)
         );
  AND2_X4 sub_436_b0_U34 ( .A1(sub_436_b0_n119), .A2(sub_436_b0_n50), .ZN(
        sub_436_b0_n34) );
  AND2_X4 sub_436_b0_U33 ( .A1(sub_436_b0_n117), .A2(sub_436_b0_n49), .ZN(
        sub_436_b0_n33) );
  AND2_X4 sub_436_b0_U32 ( .A1(sub_436_b0_n115), .A2(sub_436_b0_n48), .ZN(
        sub_436_b0_n32) );
  AND2_X4 sub_436_b0_U31 ( .A1(sub_436_b0_n113), .A2(sub_436_b0_n47), .ZN(
        sub_436_b0_n31) );
  AND2_X4 sub_436_b0_U30 ( .A1(sub_436_b0_n155), .A2(sub_436_b0_n68), .ZN(
        sub_436_b0_n30) );
  AND2_X4 sub_436_b0_U29 ( .A1(sub_436_b0_n121), .A2(sub_436_b0_n51), .ZN(
        sub_436_b0_n29) );
  AND2_X4 sub_436_b0_U28 ( .A1(sub_436_b0_n153), .A2(sub_436_b0_n67), .ZN(
        sub_436_b0_n28) );
  AND2_X4 sub_436_b0_U27 ( .A1(sub_436_b0_n109), .A2(sub_436_b0_n45), .ZN(
        sub_436_b0_n27) );
  AND2_X4 sub_436_b0_U26 ( .A1(sub_436_b0_n141), .A2(sub_436_b0_n61), .ZN(
        sub_436_b0_n26) );
  AND2_X4 sub_436_b0_U25 ( .A1(sub_436_b0_n139), .A2(sub_436_b0_n60), .ZN(
        sub_436_b0_n25) );
  AND2_X4 sub_436_b0_U24 ( .A1(sub_436_b0_n137), .A2(sub_436_b0_n59), .ZN(
        sub_436_b0_n24) );
  AND2_X4 sub_436_b0_U23 ( .A1(sub_436_b0_n135), .A2(sub_436_b0_n58), .ZN(
        sub_436_b0_n23) );
  AND2_X4 sub_436_b0_U22 ( .A1(sub_436_b0_n133), .A2(sub_436_b0_n57), .ZN(
        sub_436_b0_n22) );
  AND2_X4 sub_436_b0_U21 ( .A1(sub_436_b0_n131), .A2(sub_436_b0_n56), .ZN(
        sub_436_b0_n21) );
  AND2_X4 sub_436_b0_U20 ( .A1(sub_436_b0_n129), .A2(sub_436_b0_n55), .ZN(
        sub_436_b0_n20) );
  AND2_X4 sub_436_b0_U19 ( .A1(sub_436_b0_n127), .A2(sub_436_b0_n54), .ZN(
        sub_436_b0_n19) );
  AND2_X4 sub_436_b0_U18 ( .A1(sub_436_b0_n125), .A2(sub_436_b0_n53), .ZN(
        sub_436_b0_n18) );
  AND2_X4 sub_436_b0_U17 ( .A1(sub_436_b0_n123), .A2(sub_436_b0_n52), .ZN(
        sub_436_b0_n17) );
  AND2_X4 sub_436_b0_U16 ( .A1(sub_436_b0_n111), .A2(sub_436_b0_n46), .ZN(
        sub_436_b0_n16) );
  AND2_X4 sub_436_b0_U15 ( .A1(sub_436_b0_n151), .A2(sub_436_b0_n66), .ZN(
        sub_436_b0_n15) );
  AND2_X4 sub_436_b0_U14 ( .A1(sub_436_b0_n149), .A2(sub_436_b0_n65), .ZN(
        sub_436_b0_n14) );
  AND2_X4 sub_436_b0_U13 ( .A1(sub_436_b0_n147), .A2(sub_436_b0_n64), .ZN(
        sub_436_b0_n13) );
  AND2_X4 sub_436_b0_U12 ( .A1(sub_436_b0_n145), .A2(sub_436_b0_n63), .ZN(
        sub_436_b0_n12) );
  AND2_X4 sub_436_b0_U11 ( .A1(sub_436_b0_n143), .A2(sub_436_b0_n62), .ZN(
        sub_436_b0_n11) );
  AND2_X4 sub_436_b0_U10 ( .A1(sub_436_b0_n107), .A2(sub_436_b0_n44), .ZN(
        sub_436_b0_n10) );
  XOR2_X2 sub_436_b0_U9 ( .A(sub_436_b0_n114), .B(sub_436_b0_n32), .Z(N386) );
  XOR2_X2 sub_436_b0_U8 ( .A(sub_436_b0_n115), .B(sub_436_b0_n48), .Z(N385) );
  XOR2_X2 sub_436_b0_U7 ( .A(sub_436_b0_n116), .B(sub_436_b0_n33), .Z(N384) );
  XOR2_X2 sub_436_b0_U6 ( .A(sub_436_b0_n117), .B(sub_436_b0_n49), .Z(N383) );
  XOR2_X2 sub_436_b0_U5 ( .A(sub_436_b0_n118), .B(sub_436_b0_n34), .Z(N382) );
  XOR2_X2 sub_436_b0_U4 ( .A(sub_436_b0_n119), .B(sub_436_b0_n50), .Z(N381) );
  XOR2_X2 sub_436_b0_U3 ( .A(sub_436_b0_n120), .B(sub_436_b0_n29), .Z(N380) );
  XOR2_X2 sub_436_b0_U2 ( .A(sub_436_b0_n113), .B(sub_436_b0_n47), .Z(N387) );
  AND2_X4 sub_436_b0_U1 ( .A1(sub_436_b0_n106), .A2(sub_436_b0_n10), .ZN(
        sub_436_b0_n1) );
  AND2_X1 sll_386_U55 ( .A1(fracta_mul[0]), .A2(sll_386_n2), .ZN(
        sll_386_ML_int_1__0_) );
  AND2_X1 sll_386_U54 ( .A1(sll_386_ML_int_1__0_), .A2(sll_386_n5), .ZN(
        sll_386_ML_int_2__0_) );
  AND2_X1 sll_386_U53 ( .A1(sll_386_ML_int_1__1_), .A2(sll_386_n5), .ZN(
        sll_386_ML_int_2__1_) );
  AND2_X1 sll_386_U52 ( .A1(sll_386_ML_int_2__0_), .A2(sll_386_n8), .ZN(
        sll_386_ML_int_3__0_) );
  AND2_X1 sll_386_U51 ( .A1(sll_386_ML_int_2__1_), .A2(sll_386_n8), .ZN(
        sll_386_ML_int_3__1_) );
  AND2_X1 sll_386_U50 ( .A1(sll_386_ML_int_2__2_), .A2(sll_386_n8), .ZN(
        sll_386_ML_int_3__2_) );
  AND2_X1 sll_386_U49 ( .A1(sll_386_ML_int_2__3_), .A2(sll_386_n8), .ZN(
        sll_386_ML_int_3__3_) );
  NAND2_X1 sll_386_U48 ( .A1(sll_386_ML_int_3__0_), .A2(sll_386_n10), .ZN(
        sll_386_n30) );
  NAND2_X1 sll_386_U47 ( .A1(sll_386_ML_int_3__1_), .A2(sll_386_n10), .ZN(
        sll_386_n29) );
  NAND2_X1 sll_386_U46 ( .A1(sll_386_ML_int_3__2_), .A2(sll_386_n10), .ZN(
        sll_386_n28) );
  NAND2_X1 sll_386_U45 ( .A1(sll_386_ML_int_3__3_), .A2(sll_386_n10), .ZN(
        sll_386_n27) );
  NAND2_X1 sll_386_U44 ( .A1(sll_386_ML_int_3__4_), .A2(sll_386_n10), .ZN(
        sll_386_n26) );
  NAND2_X1 sll_386_U43 ( .A1(sll_386_ML_int_3__5_), .A2(sll_386_n10), .ZN(
        sll_386_n25) );
  NAND2_X1 sll_386_U42 ( .A1(sll_386_ML_int_3__6_), .A2(sll_386_n10), .ZN(
        sll_386_n24) );
  NAND2_X1 sll_386_U41 ( .A1(sll_386_ML_int_3__7_), .A2(sll_386_n10), .ZN(
        sll_386_n23) );
  NOR2_X1 sll_386_U40 ( .A1(div_opa_ldz_d[4]), .A2(sll_386_n30), .ZN(N256) );
  AND2_X1 sll_386_U39 ( .A1(sll_386_ML_int_4__10_), .A2(sll_386_n12), .ZN(N266) );
  AND2_X1 sll_386_U38 ( .A1(sll_386_ML_int_4__11_), .A2(sll_386_n12), .ZN(N267) );
  AND2_X1 sll_386_U37 ( .A1(sll_386_ML_int_4__12_), .A2(sll_386_n12), .ZN(N268) );
  AND2_X1 sll_386_U36 ( .A1(sll_386_ML_int_4__13_), .A2(sll_386_n12), .ZN(N269) );
  AND2_X1 sll_386_U35 ( .A1(sll_386_ML_int_4__14_), .A2(sll_386_n12), .ZN(N270) );
  AND2_X1 sll_386_U34 ( .A1(sll_386_ML_int_4__15_), .A2(sll_386_n12), .ZN(N271) );
  NOR2_X1 sll_386_U33 ( .A1(sll_386_n13), .A2(sll_386_n29), .ZN(N257) );
  NOR2_X1 sll_386_U32 ( .A1(sll_386_n14), .A2(sll_386_n28), .ZN(N258) );
  NOR2_X1 sll_386_U31 ( .A1(sll_386_n11), .A2(sll_386_n27), .ZN(N259) );
  NOR2_X1 sll_386_U30 ( .A1(sll_386_n11), .A2(sll_386_n26), .ZN(N260) );
  NOR2_X1 sll_386_U29 ( .A1(sll_386_n11), .A2(sll_386_n25), .ZN(N261) );
  NOR2_X1 sll_386_U28 ( .A1(sll_386_n11), .A2(sll_386_n24), .ZN(N262) );
  NOR2_X1 sll_386_U27 ( .A1(sll_386_n11), .A2(sll_386_n23), .ZN(N263) );
  AND2_X1 sll_386_U26 ( .A1(sll_386_ML_int_4__8_), .A2(sll_386_n12), .ZN(N264)
         );
  AND2_X1 sll_386_U25 ( .A1(sll_386_ML_int_4__9_), .A2(sll_386_n12), .ZN(N265)
         );
  INV_X4 sll_386_U24 ( .A(sll_386_n23), .ZN(sll_386_n22) );
  INV_X4 sll_386_U23 ( .A(sll_386_n24), .ZN(sll_386_n21) );
  INV_X4 sll_386_U22 ( .A(sll_386_n25), .ZN(sll_386_n20) );
  INV_X4 sll_386_U21 ( .A(sll_386_n26), .ZN(sll_386_n19) );
  INV_X4 sll_386_U20 ( .A(sll_386_n30), .ZN(sll_386_n18) );
  INV_X4 sll_386_U19 ( .A(sll_386_n29), .ZN(sll_386_n17) );
  INV_X4 sll_386_U18 ( .A(sll_386_n28), .ZN(sll_386_n16) );
  INV_X4 sll_386_U17 ( .A(sll_386_n27), .ZN(sll_386_n15) );
  INV_X4 sll_386_U16 ( .A(sll_386_n10), .ZN(sll_386_n9) );
  INV_X4 sll_386_U15 ( .A(sll_386_n12), .ZN(sll_386_n13) );
  INV_X4 sll_386_U14 ( .A(sll_386_n12), .ZN(sll_386_n14) );
  INV_X4 sll_386_U13 ( .A(sll_386_n12), .ZN(sll_386_n11) );
  INV_X4 sll_386_U12 ( .A(sll_386_n8), .ZN(sll_386_n7) );
  INV_X4 sll_386_U11 ( .A(div_opa_ldz_d[1]), .ZN(sll_386_n5) );
  INV_X4 sll_386_U10 ( .A(sll_386_n5), .ZN(sll_386_n4) );
  INV_X4 sll_386_U9 ( .A(div_opa_ldz_d[0]), .ZN(sll_386_n2) );
  INV_X4 sll_386_U8 ( .A(sll_386_n2), .ZN(sll_386_n1) );
  INV_X4 sll_386_U7 ( .A(div_opa_ldz_d[4]), .ZN(sll_386_n12) );
  INV_X4 sll_386_U6 ( .A(sll_386_n2), .ZN(sll_386_n3) );
  INV_X4 sll_386_U5 ( .A(sll_386_n5), .ZN(sll_386_n6) );
  INV_X4 sll_386_U4 ( .A(div_opa_ldz_d[2]), .ZN(sll_386_n8) );
  INV_X4 sll_386_U3 ( .A(div_opa_ldz_d[3]), .ZN(sll_386_n10) );
  MUX2_X2 sll_386_M1_0_1 ( .A(fracta_mul[1]), .B(fracta_mul[0]), .S(sll_386_n3), .Z(sll_386_ML_int_1__1_) );
  MUX2_X2 sll_386_M1_0_2 ( .A(fracta_mul[2]), .B(fracta_mul[1]), .S(sll_386_n3), .Z(sll_386_ML_int_1__2_) );
  MUX2_X2 sll_386_M1_0_3 ( .A(fracta_mul[3]), .B(fracta_mul[2]), .S(sll_386_n3), .Z(sll_386_ML_int_1__3_) );
  MUX2_X2 sll_386_M1_0_4 ( .A(fracta_mul[4]), .B(fracta_mul[3]), .S(sll_386_n3), .Z(sll_386_ML_int_1__4_) );
  MUX2_X2 sll_386_M1_0_5 ( .A(fracta_mul[5]), .B(fracta_mul[4]), .S(sll_386_n3), .Z(sll_386_ML_int_1__5_) );
  MUX2_X2 sll_386_M1_0_6 ( .A(fracta_mul[6]), .B(fracta_mul[5]), .S(sll_386_n3), .Z(sll_386_ML_int_1__6_) );
  MUX2_X2 sll_386_M1_0_7 ( .A(fracta_mul[7]), .B(fracta_mul[6]), .S(sll_386_n3), .Z(sll_386_ML_int_1__7_) );
  MUX2_X2 sll_386_M1_0_8 ( .A(fracta_mul[8]), .B(fracta_mul[7]), .S(sll_386_n3), .Z(sll_386_ML_int_1__8_) );
  MUX2_X2 sll_386_M1_0_9 ( .A(fracta_mul[9]), .B(fracta_mul[8]), .S(sll_386_n3), .Z(sll_386_ML_int_1__9_) );
  MUX2_X2 sll_386_M1_0_10 ( .A(fracta_mul[10]), .B(fracta_mul[9]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__10_) );
  MUX2_X2 sll_386_M1_0_11 ( .A(fracta_mul[11]), .B(fracta_mul[10]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__11_) );
  MUX2_X2 sll_386_M1_0_12 ( .A(fracta_mul[12]), .B(fracta_mul[11]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__12_) );
  MUX2_X2 sll_386_M1_0_13 ( .A(fracta_mul[13]), .B(fracta_mul[12]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__13_) );
  MUX2_X2 sll_386_M1_0_14 ( .A(fracta_mul[14]), .B(fracta_mul[13]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__14_) );
  MUX2_X2 sll_386_M1_0_15 ( .A(fracta_mul[15]), .B(fracta_mul[14]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__15_) );
  MUX2_X2 sll_386_M1_0_16 ( .A(fracta_mul[16]), .B(fracta_mul[15]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__16_) );
  MUX2_X2 sll_386_M1_0_17 ( .A(fracta_mul[17]), .B(fracta_mul[16]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__17_) );
  MUX2_X2 sll_386_M1_0_18 ( .A(fracta_mul[18]), .B(fracta_mul[17]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__18_) );
  MUX2_X2 sll_386_M1_0_19 ( .A(fracta_mul[19]), .B(fracta_mul[18]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__19_) );
  MUX2_X2 sll_386_M1_0_20 ( .A(fracta_mul[20]), .B(fracta_mul[19]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__20_) );
  MUX2_X2 sll_386_M1_0_21 ( .A(fracta_mul[21]), .B(fracta_mul[20]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__21_) );
  MUX2_X2 sll_386_M1_0_22 ( .A(fracta_mul[22]), .B(fracta_mul[21]), .S(
        sll_386_n3), .Z(sll_386_ML_int_1__22_) );
  MUX2_X2 sll_386_M1_0_23 ( .A(fracta_mul[23]), .B(fracta_mul[22]), .S(
        div_opa_ldz_d[0]), .Z(sll_386_ML_int_1__23_) );
  MUX2_X2 sll_386_M1_0_24 ( .A(fracta_mul[24]), .B(fracta_mul[23]), .S(
        div_opa_ldz_d[0]), .Z(sll_386_ML_int_1__24_) );
  MUX2_X2 sll_386_M1_0_25 ( .A(fracta_mul[25]), .B(fracta_mul[24]), .S(
        sll_386_n1), .Z(sll_386_ML_int_1__25_) );
  MUX2_X2 sll_386_M1_0_26 ( .A(fracta_mul[26]), .B(fracta_mul[25]), .S(
        sll_386_n1), .Z(sll_386_ML_int_1__26_) );
  MUX2_X2 sll_386_M1_0_27 ( .A(fracta_mul[27]), .B(fracta_mul[26]), .S(
        div_opa_ldz_d[0]), .Z(sll_386_ML_int_1__27_) );
  MUX2_X2 sll_386_M1_0_28 ( .A(fracta_mul[28]), .B(fracta_mul[27]), .S(
        div_opa_ldz_d[0]), .Z(sll_386_ML_int_1__28_) );
  MUX2_X2 sll_386_M1_0_29 ( .A(fracta_mul[29]), .B(fracta_mul[28]), .S(
        div_opa_ldz_d[0]), .Z(sll_386_ML_int_1__29_) );
  MUX2_X2 sll_386_M1_0_30 ( .A(fracta_mul[30]), .B(fracta_mul[29]), .S(
        div_opa_ldz_d[0]), .Z(sll_386_ML_int_1__30_) );
  MUX2_X2 sll_386_M1_0_31 ( .A(fracta_mul[31]), .B(fracta_mul[30]), .S(
        div_opa_ldz_d[0]), .Z(sll_386_ML_int_1__31_) );
  MUX2_X2 sll_386_M1_0_32 ( .A(fracta_mul[32]), .B(fracta_mul[31]), .S(
        div_opa_ldz_d[0]), .Z(sll_386_ML_int_1__32_) );
  MUX2_X2 sll_386_M1_0_33 ( .A(fracta_mul[33]), .B(fracta_mul[32]), .S(
        div_opa_ldz_d[0]), .Z(sll_386_ML_int_1__33_) );
  MUX2_X2 sll_386_M1_0_34 ( .A(fracta_mul[34]), .B(fracta_mul[33]), .S(
        div_opa_ldz_d[0]), .Z(sll_386_ML_int_1__34_) );
  MUX2_X2 sll_386_M1_0_35 ( .A(fracta_mul[35]), .B(fracta_mul[34]), .S(
        div_opa_ldz_d[0]), .Z(sll_386_ML_int_1__35_) );
  MUX2_X2 sll_386_M1_0_36 ( .A(fracta_mul[36]), .B(fracta_mul[35]), .S(
        div_opa_ldz_d[0]), .Z(sll_386_ML_int_1__36_) );
  MUX2_X2 sll_386_M1_0_37 ( .A(fracta_mul[37]), .B(fracta_mul[36]), .S(
        div_opa_ldz_d[0]), .Z(sll_386_ML_int_1__37_) );
  MUX2_X2 sll_386_M1_0_38 ( .A(fracta_mul[38]), .B(fracta_mul[37]), .S(
        div_opa_ldz_d[0]), .Z(sll_386_ML_int_1__38_) );
  MUX2_X2 sll_386_M1_0_39 ( .A(fracta_mul[39]), .B(fracta_mul[38]), .S(
        div_opa_ldz_d[0]), .Z(sll_386_ML_int_1__39_) );
  MUX2_X2 sll_386_M1_0_40 ( .A(fracta_mul[40]), .B(fracta_mul[39]), .S(
        div_opa_ldz_d[0]), .Z(sll_386_ML_int_1__40_) );
  MUX2_X2 sll_386_M1_0_41 ( .A(fracta_mul[41]), .B(fracta_mul[40]), .S(
        div_opa_ldz_d[0]), .Z(sll_386_ML_int_1__41_) );
  MUX2_X2 sll_386_M1_0_42 ( .A(fracta_mul[42]), .B(fracta_mul[41]), .S(
        div_opa_ldz_d[0]), .Z(sll_386_ML_int_1__42_) );
  MUX2_X2 sll_386_M1_0_43 ( .A(fracta_mul[43]), .B(fracta_mul[42]), .S(
        div_opa_ldz_d[0]), .Z(sll_386_ML_int_1__43_) );
  MUX2_X2 sll_386_M1_0_44 ( .A(fracta_mul[44]), .B(fracta_mul[43]), .S(
        div_opa_ldz_d[0]), .Z(sll_386_ML_int_1__44_) );
  MUX2_X2 sll_386_M1_0_45 ( .A(fracta_mul[45]), .B(fracta_mul[44]), .S(
        div_opa_ldz_d[0]), .Z(sll_386_ML_int_1__45_) );
  MUX2_X2 sll_386_M1_0_46 ( .A(fracta_mul[46]), .B(fracta_mul[45]), .S(
        div_opa_ldz_d[0]), .Z(sll_386_ML_int_1__46_) );
  MUX2_X2 sll_386_M1_0_47 ( .A(fracta_mul[47]), .B(fracta_mul[46]), .S(
        div_opa_ldz_d[0]), .Z(sll_386_ML_int_1__47_) );
  MUX2_X2 sll_386_M1_0_48 ( .A(fracta_mul[48]), .B(fracta_mul[47]), .S(
        sll_386_n1), .Z(sll_386_ML_int_1__48_) );
  MUX2_X2 sll_386_M1_0_49 ( .A(fracta_mul[49]), .B(fracta_mul[48]), .S(
        sll_386_n1), .Z(sll_386_ML_int_1__49_) );
  MUX2_X2 sll_386_M1_0_50 ( .A(fracta_mul[50]), .B(fracta_mul[49]), .S(
        sll_386_n1), .Z(sll_386_ML_int_1__50_) );
  MUX2_X2 sll_386_M1_0_51 ( .A(fracta_mul[51]), .B(fracta_mul[50]), .S(
        sll_386_n1), .Z(sll_386_ML_int_1__51_) );
  MUX2_X2 sll_386_M1_0_52 ( .A(n4602), .B(fracta_mul[51]), .S(sll_386_n1), .Z(
        sll_386_ML_int_1__52_) );
  MUX2_X2 sll_386_M1_1_2 ( .A(sll_386_ML_int_1__2_), .B(sll_386_ML_int_1__0_), 
        .S(sll_386_n6), .Z(sll_386_ML_int_2__2_) );
  MUX2_X2 sll_386_M1_1_3 ( .A(sll_386_ML_int_1__3_), .B(sll_386_ML_int_1__1_), 
        .S(sll_386_n6), .Z(sll_386_ML_int_2__3_) );
  MUX2_X2 sll_386_M1_1_4 ( .A(sll_386_ML_int_1__4_), .B(sll_386_ML_int_1__2_), 
        .S(sll_386_n6), .Z(sll_386_ML_int_2__4_) );
  MUX2_X2 sll_386_M1_1_5 ( .A(sll_386_ML_int_1__5_), .B(sll_386_ML_int_1__3_), 
        .S(sll_386_n6), .Z(sll_386_ML_int_2__5_) );
  MUX2_X2 sll_386_M1_1_6 ( .A(sll_386_ML_int_1__6_), .B(sll_386_ML_int_1__4_), 
        .S(sll_386_n6), .Z(sll_386_ML_int_2__6_) );
  MUX2_X2 sll_386_M1_1_7 ( .A(sll_386_ML_int_1__7_), .B(sll_386_ML_int_1__5_), 
        .S(sll_386_n6), .Z(sll_386_ML_int_2__7_) );
  MUX2_X2 sll_386_M1_1_8 ( .A(sll_386_ML_int_1__8_), .B(sll_386_ML_int_1__6_), 
        .S(sll_386_n6), .Z(sll_386_ML_int_2__8_) );
  MUX2_X2 sll_386_M1_1_9 ( .A(sll_386_ML_int_1__9_), .B(sll_386_ML_int_1__7_), 
        .S(sll_386_n6), .Z(sll_386_ML_int_2__9_) );
  MUX2_X2 sll_386_M1_1_10 ( .A(sll_386_ML_int_1__10_), .B(sll_386_ML_int_1__8_), .S(sll_386_n6), .Z(sll_386_ML_int_2__10_) );
  MUX2_X2 sll_386_M1_1_11 ( .A(sll_386_ML_int_1__11_), .B(sll_386_ML_int_1__9_), .S(sll_386_n6), .Z(sll_386_ML_int_2__11_) );
  MUX2_X2 sll_386_M1_1_12 ( .A(sll_386_ML_int_1__12_), .B(
        sll_386_ML_int_1__10_), .S(sll_386_n6), .Z(sll_386_ML_int_2__12_) );
  MUX2_X2 sll_386_M1_1_13 ( .A(sll_386_ML_int_1__13_), .B(
        sll_386_ML_int_1__11_), .S(sll_386_n6), .Z(sll_386_ML_int_2__13_) );
  MUX2_X2 sll_386_M1_1_14 ( .A(sll_386_ML_int_1__14_), .B(
        sll_386_ML_int_1__12_), .S(sll_386_n6), .Z(sll_386_ML_int_2__14_) );
  MUX2_X2 sll_386_M1_1_15 ( .A(sll_386_ML_int_1__15_), .B(
        sll_386_ML_int_1__13_), .S(sll_386_n6), .Z(sll_386_ML_int_2__15_) );
  MUX2_X2 sll_386_M1_1_16 ( .A(sll_386_ML_int_1__16_), .B(
        sll_386_ML_int_1__14_), .S(sll_386_n6), .Z(sll_386_ML_int_2__16_) );
  MUX2_X2 sll_386_M1_1_17 ( .A(sll_386_ML_int_1__17_), .B(
        sll_386_ML_int_1__15_), .S(sll_386_n6), .Z(sll_386_ML_int_2__17_) );
  MUX2_X2 sll_386_M1_1_18 ( .A(sll_386_ML_int_1__18_), .B(
        sll_386_ML_int_1__16_), .S(sll_386_n6), .Z(sll_386_ML_int_2__18_) );
  MUX2_X2 sll_386_M1_1_19 ( .A(sll_386_ML_int_1__19_), .B(
        sll_386_ML_int_1__17_), .S(sll_386_n6), .Z(sll_386_ML_int_2__19_) );
  MUX2_X2 sll_386_M1_1_20 ( .A(sll_386_ML_int_1__20_), .B(
        sll_386_ML_int_1__18_), .S(sll_386_n6), .Z(sll_386_ML_int_2__20_) );
  MUX2_X2 sll_386_M1_1_21 ( .A(sll_386_ML_int_1__21_), .B(
        sll_386_ML_int_1__19_), .S(sll_386_n6), .Z(sll_386_ML_int_2__21_) );
  MUX2_X2 sll_386_M1_1_22 ( .A(sll_386_ML_int_1__22_), .B(
        sll_386_ML_int_1__20_), .S(sll_386_n6), .Z(sll_386_ML_int_2__22_) );
  MUX2_X2 sll_386_M1_1_23 ( .A(sll_386_ML_int_1__23_), .B(
        sll_386_ML_int_1__21_), .S(sll_386_n6), .Z(sll_386_ML_int_2__23_) );
  MUX2_X2 sll_386_M1_1_24 ( .A(sll_386_ML_int_1__24_), .B(
        sll_386_ML_int_1__22_), .S(div_opa_ldz_d[1]), .Z(sll_386_ML_int_2__24_) );
  MUX2_X2 sll_386_M1_1_25 ( .A(sll_386_ML_int_1__25_), .B(
        sll_386_ML_int_1__23_), .S(div_opa_ldz_d[1]), .Z(sll_386_ML_int_2__25_) );
  MUX2_X2 sll_386_M1_1_26 ( .A(sll_386_ML_int_1__26_), .B(
        sll_386_ML_int_1__24_), .S(div_opa_ldz_d[1]), .Z(sll_386_ML_int_2__26_) );
  MUX2_X2 sll_386_M1_1_27 ( .A(sll_386_ML_int_1__27_), .B(
        sll_386_ML_int_1__25_), .S(sll_386_n4), .Z(sll_386_ML_int_2__27_) );
  MUX2_X2 sll_386_M1_1_28 ( .A(sll_386_ML_int_1__28_), .B(
        sll_386_ML_int_1__26_), .S(sll_386_n4), .Z(sll_386_ML_int_2__28_) );
  MUX2_X2 sll_386_M1_1_29 ( .A(sll_386_ML_int_1__29_), .B(
        sll_386_ML_int_1__27_), .S(div_opa_ldz_d[1]), .Z(sll_386_ML_int_2__29_) );
  MUX2_X2 sll_386_M1_1_30 ( .A(sll_386_ML_int_1__30_), .B(
        sll_386_ML_int_1__28_), .S(div_opa_ldz_d[1]), .Z(sll_386_ML_int_2__30_) );
  MUX2_X2 sll_386_M1_1_31 ( .A(sll_386_ML_int_1__31_), .B(
        sll_386_ML_int_1__29_), .S(div_opa_ldz_d[1]), .Z(sll_386_ML_int_2__31_) );
  MUX2_X2 sll_386_M1_1_32 ( .A(sll_386_ML_int_1__32_), .B(
        sll_386_ML_int_1__30_), .S(div_opa_ldz_d[1]), .Z(sll_386_ML_int_2__32_) );
  MUX2_X2 sll_386_M1_1_33 ( .A(sll_386_ML_int_1__33_), .B(
        sll_386_ML_int_1__31_), .S(div_opa_ldz_d[1]), .Z(sll_386_ML_int_2__33_) );
  MUX2_X2 sll_386_M1_1_34 ( .A(sll_386_ML_int_1__34_), .B(
        sll_386_ML_int_1__32_), .S(div_opa_ldz_d[1]), .Z(sll_386_ML_int_2__34_) );
  MUX2_X2 sll_386_M1_1_35 ( .A(sll_386_ML_int_1__35_), .B(
        sll_386_ML_int_1__33_), .S(div_opa_ldz_d[1]), .Z(sll_386_ML_int_2__35_) );
  MUX2_X2 sll_386_M1_1_36 ( .A(sll_386_ML_int_1__36_), .B(
        sll_386_ML_int_1__34_), .S(div_opa_ldz_d[1]), .Z(sll_386_ML_int_2__36_) );
  MUX2_X2 sll_386_M1_1_37 ( .A(sll_386_ML_int_1__37_), .B(
        sll_386_ML_int_1__35_), .S(div_opa_ldz_d[1]), .Z(sll_386_ML_int_2__37_) );
  MUX2_X2 sll_386_M1_1_38 ( .A(sll_386_ML_int_1__38_), .B(
        sll_386_ML_int_1__36_), .S(div_opa_ldz_d[1]), .Z(sll_386_ML_int_2__38_) );
  MUX2_X2 sll_386_M1_1_39 ( .A(sll_386_ML_int_1__39_), .B(
        sll_386_ML_int_1__37_), .S(div_opa_ldz_d[1]), .Z(sll_386_ML_int_2__39_) );
  MUX2_X2 sll_386_M1_1_40 ( .A(sll_386_ML_int_1__40_), .B(
        sll_386_ML_int_1__38_), .S(div_opa_ldz_d[1]), .Z(sll_386_ML_int_2__40_) );
  MUX2_X2 sll_386_M1_1_41 ( .A(sll_386_ML_int_1__41_), .B(
        sll_386_ML_int_1__39_), .S(div_opa_ldz_d[1]), .Z(sll_386_ML_int_2__41_) );
  MUX2_X2 sll_386_M1_1_42 ( .A(sll_386_ML_int_1__42_), .B(
        sll_386_ML_int_1__40_), .S(div_opa_ldz_d[1]), .Z(sll_386_ML_int_2__42_) );
  MUX2_X2 sll_386_M1_1_43 ( .A(sll_386_ML_int_1__43_), .B(
        sll_386_ML_int_1__41_), .S(div_opa_ldz_d[1]), .Z(sll_386_ML_int_2__43_) );
  MUX2_X2 sll_386_M1_1_44 ( .A(sll_386_ML_int_1__44_), .B(
        sll_386_ML_int_1__42_), .S(div_opa_ldz_d[1]), .Z(sll_386_ML_int_2__44_) );
  MUX2_X2 sll_386_M1_1_45 ( .A(sll_386_ML_int_1__45_), .B(
        sll_386_ML_int_1__43_), .S(div_opa_ldz_d[1]), .Z(sll_386_ML_int_2__45_) );
  MUX2_X2 sll_386_M1_1_46 ( .A(sll_386_ML_int_1__46_), .B(
        sll_386_ML_int_1__44_), .S(div_opa_ldz_d[1]), .Z(sll_386_ML_int_2__46_) );
  MUX2_X2 sll_386_M1_1_47 ( .A(sll_386_ML_int_1__47_), .B(
        sll_386_ML_int_1__45_), .S(div_opa_ldz_d[1]), .Z(sll_386_ML_int_2__47_) );
  MUX2_X2 sll_386_M1_1_48 ( .A(sll_386_ML_int_1__48_), .B(
        sll_386_ML_int_1__46_), .S(div_opa_ldz_d[1]), .Z(sll_386_ML_int_2__48_) );
  MUX2_X2 sll_386_M1_1_49 ( .A(sll_386_ML_int_1__49_), .B(
        sll_386_ML_int_1__47_), .S(sll_386_n4), .Z(sll_386_ML_int_2__49_) );
  MUX2_X2 sll_386_M1_1_50 ( .A(sll_386_ML_int_1__50_), .B(
        sll_386_ML_int_1__48_), .S(sll_386_n4), .Z(sll_386_ML_int_2__50_) );
  MUX2_X2 sll_386_M1_1_51 ( .A(sll_386_ML_int_1__51_), .B(
        sll_386_ML_int_1__49_), .S(sll_386_n4), .Z(sll_386_ML_int_2__51_) );
  MUX2_X2 sll_386_M1_1_52 ( .A(sll_386_ML_int_1__52_), .B(
        sll_386_ML_int_1__50_), .S(sll_386_n4), .Z(sll_386_ML_int_2__52_) );
  MUX2_X2 sll_386_M1_2_4 ( .A(sll_386_ML_int_2__4_), .B(sll_386_ML_int_2__0_), 
        .S(div_opa_ldz_d[2]), .Z(sll_386_ML_int_3__4_) );
  MUX2_X2 sll_386_M1_2_5 ( .A(sll_386_ML_int_2__5_), .B(sll_386_ML_int_2__1_), 
        .S(div_opa_ldz_d[2]), .Z(sll_386_ML_int_3__5_) );
  MUX2_X2 sll_386_M1_2_6 ( .A(sll_386_ML_int_2__6_), .B(sll_386_ML_int_2__2_), 
        .S(div_opa_ldz_d[2]), .Z(sll_386_ML_int_3__6_) );
  MUX2_X2 sll_386_M1_2_7 ( .A(sll_386_ML_int_2__7_), .B(sll_386_ML_int_2__3_), 
        .S(div_opa_ldz_d[2]), .Z(sll_386_ML_int_3__7_) );
  MUX2_X2 sll_386_M1_2_8 ( .A(sll_386_ML_int_2__8_), .B(sll_386_ML_int_2__4_), 
        .S(div_opa_ldz_d[2]), .Z(sll_386_ML_int_3__8_) );
  MUX2_X2 sll_386_M1_2_9 ( .A(sll_386_ML_int_2__9_), .B(sll_386_ML_int_2__5_), 
        .S(div_opa_ldz_d[2]), .Z(sll_386_ML_int_3__9_) );
  MUX2_X2 sll_386_M1_2_10 ( .A(sll_386_ML_int_2__10_), .B(sll_386_ML_int_2__6_), .S(div_opa_ldz_d[2]), .Z(sll_386_ML_int_3__10_) );
  MUX2_X2 sll_386_M1_2_11 ( .A(sll_386_ML_int_2__11_), .B(sll_386_ML_int_2__7_), .S(div_opa_ldz_d[2]), .Z(sll_386_ML_int_3__11_) );
  MUX2_X2 sll_386_M1_2_12 ( .A(sll_386_ML_int_2__12_), .B(sll_386_ML_int_2__8_), .S(div_opa_ldz_d[2]), .Z(sll_386_ML_int_3__12_) );
  MUX2_X2 sll_386_M1_2_13 ( .A(sll_386_ML_int_2__13_), .B(sll_386_ML_int_2__9_), .S(div_opa_ldz_d[2]), .Z(sll_386_ML_int_3__13_) );
  MUX2_X2 sll_386_M1_2_14 ( .A(sll_386_ML_int_2__14_), .B(
        sll_386_ML_int_2__10_), .S(div_opa_ldz_d[2]), .Z(sll_386_ML_int_3__14_) );
  MUX2_X2 sll_386_M1_2_15 ( .A(sll_386_ML_int_2__15_), .B(
        sll_386_ML_int_2__11_), .S(div_opa_ldz_d[2]), .Z(sll_386_ML_int_3__15_) );
  MUX2_X2 sll_386_M1_2_16 ( .A(sll_386_ML_int_2__16_), .B(
        sll_386_ML_int_2__12_), .S(div_opa_ldz_d[2]), .Z(sll_386_ML_int_3__16_) );
  MUX2_X2 sll_386_M1_2_17 ( .A(sll_386_ML_int_2__17_), .B(
        sll_386_ML_int_2__13_), .S(div_opa_ldz_d[2]), .Z(sll_386_ML_int_3__17_) );
  MUX2_X2 sll_386_M1_2_18 ( .A(sll_386_ML_int_2__18_), .B(
        sll_386_ML_int_2__14_), .S(div_opa_ldz_d[2]), .Z(sll_386_ML_int_3__18_) );
  MUX2_X2 sll_386_M1_2_19 ( .A(sll_386_ML_int_2__19_), .B(
        sll_386_ML_int_2__15_), .S(div_opa_ldz_d[2]), .Z(sll_386_ML_int_3__19_) );
  MUX2_X2 sll_386_M1_2_20 ( .A(sll_386_ML_int_2__20_), .B(
        sll_386_ML_int_2__16_), .S(div_opa_ldz_d[2]), .Z(sll_386_ML_int_3__20_) );
  MUX2_X2 sll_386_M1_2_21 ( .A(sll_386_ML_int_2__21_), .B(
        sll_386_ML_int_2__17_), .S(div_opa_ldz_d[2]), .Z(sll_386_ML_int_3__21_) );
  MUX2_X2 sll_386_M1_2_22 ( .A(sll_386_ML_int_2__22_), .B(
        sll_386_ML_int_2__18_), .S(div_opa_ldz_d[2]), .Z(sll_386_ML_int_3__22_) );
  MUX2_X2 sll_386_M1_2_23 ( .A(sll_386_ML_int_2__23_), .B(
        sll_386_ML_int_2__19_), .S(div_opa_ldz_d[2]), .Z(sll_386_ML_int_3__23_) );
  MUX2_X2 sll_386_M1_2_24 ( .A(sll_386_ML_int_2__24_), .B(
        sll_386_ML_int_2__20_), .S(div_opa_ldz_d[2]), .Z(sll_386_ML_int_3__24_) );
  MUX2_X2 sll_386_M1_2_25 ( .A(sll_386_ML_int_2__25_), .B(
        sll_386_ML_int_2__21_), .S(div_opa_ldz_d[2]), .Z(sll_386_ML_int_3__25_) );
  MUX2_X2 sll_386_M1_2_26 ( .A(sll_386_ML_int_2__26_), .B(
        sll_386_ML_int_2__22_), .S(sll_386_n7), .Z(sll_386_ML_int_3__26_) );
  MUX2_X2 sll_386_M1_2_27 ( .A(sll_386_ML_int_2__27_), .B(
        sll_386_ML_int_2__23_), .S(sll_386_n7), .Z(sll_386_ML_int_3__27_) );
  MUX2_X2 sll_386_M1_2_28 ( .A(sll_386_ML_int_2__28_), .B(
        sll_386_ML_int_2__24_), .S(sll_386_n7), .Z(sll_386_ML_int_3__28_) );
  MUX2_X2 sll_386_M1_2_29 ( .A(sll_386_ML_int_2__29_), .B(
        sll_386_ML_int_2__25_), .S(sll_386_n7), .Z(sll_386_ML_int_3__29_) );
  MUX2_X2 sll_386_M1_2_30 ( .A(sll_386_ML_int_2__30_), .B(
        sll_386_ML_int_2__26_), .S(sll_386_n7), .Z(sll_386_ML_int_3__30_) );
  MUX2_X2 sll_386_M1_2_31 ( .A(sll_386_ML_int_2__31_), .B(
        sll_386_ML_int_2__27_), .S(sll_386_n7), .Z(sll_386_ML_int_3__31_) );
  MUX2_X2 sll_386_M1_2_32 ( .A(sll_386_ML_int_2__32_), .B(
        sll_386_ML_int_2__28_), .S(sll_386_n7), .Z(sll_386_ML_int_3__32_) );
  MUX2_X2 sll_386_M1_2_33 ( .A(sll_386_ML_int_2__33_), .B(
        sll_386_ML_int_2__29_), .S(sll_386_n7), .Z(sll_386_ML_int_3__33_) );
  MUX2_X2 sll_386_M1_2_34 ( .A(sll_386_ML_int_2__34_), .B(
        sll_386_ML_int_2__30_), .S(sll_386_n7), .Z(sll_386_ML_int_3__34_) );
  MUX2_X2 sll_386_M1_2_35 ( .A(sll_386_ML_int_2__35_), .B(
        sll_386_ML_int_2__31_), .S(sll_386_n7), .Z(sll_386_ML_int_3__35_) );
  MUX2_X2 sll_386_M1_2_36 ( .A(sll_386_ML_int_2__36_), .B(
        sll_386_ML_int_2__32_), .S(sll_386_n7), .Z(sll_386_ML_int_3__36_) );
  MUX2_X2 sll_386_M1_2_37 ( .A(sll_386_ML_int_2__37_), .B(
        sll_386_ML_int_2__33_), .S(sll_386_n7), .Z(sll_386_ML_int_3__37_) );
  MUX2_X2 sll_386_M1_2_38 ( .A(sll_386_ML_int_2__38_), .B(
        sll_386_ML_int_2__34_), .S(sll_386_n7), .Z(sll_386_ML_int_3__38_) );
  MUX2_X2 sll_386_M1_2_39 ( .A(sll_386_ML_int_2__39_), .B(
        sll_386_ML_int_2__35_), .S(sll_386_n7), .Z(sll_386_ML_int_3__39_) );
  MUX2_X2 sll_386_M1_2_40 ( .A(sll_386_ML_int_2__40_), .B(
        sll_386_ML_int_2__36_), .S(sll_386_n7), .Z(sll_386_ML_int_3__40_) );
  MUX2_X2 sll_386_M1_2_41 ( .A(sll_386_ML_int_2__41_), .B(
        sll_386_ML_int_2__37_), .S(sll_386_n7), .Z(sll_386_ML_int_3__41_) );
  MUX2_X2 sll_386_M1_2_42 ( .A(sll_386_ML_int_2__42_), .B(
        sll_386_ML_int_2__38_), .S(sll_386_n7), .Z(sll_386_ML_int_3__42_) );
  MUX2_X2 sll_386_M1_2_43 ( .A(sll_386_ML_int_2__43_), .B(
        sll_386_ML_int_2__39_), .S(sll_386_n7), .Z(sll_386_ML_int_3__43_) );
  MUX2_X2 sll_386_M1_2_44 ( .A(sll_386_ML_int_2__44_), .B(
        sll_386_ML_int_2__40_), .S(sll_386_n7), .Z(sll_386_ML_int_3__44_) );
  MUX2_X2 sll_386_M1_2_45 ( .A(sll_386_ML_int_2__45_), .B(
        sll_386_ML_int_2__41_), .S(sll_386_n7), .Z(sll_386_ML_int_3__45_) );
  MUX2_X2 sll_386_M1_2_46 ( .A(sll_386_ML_int_2__46_), .B(
        sll_386_ML_int_2__42_), .S(sll_386_n7), .Z(sll_386_ML_int_3__46_) );
  MUX2_X2 sll_386_M1_2_47 ( .A(sll_386_ML_int_2__47_), .B(
        sll_386_ML_int_2__43_), .S(sll_386_n7), .Z(sll_386_ML_int_3__47_) );
  MUX2_X2 sll_386_M1_2_48 ( .A(sll_386_ML_int_2__48_), .B(
        sll_386_ML_int_2__44_), .S(sll_386_n7), .Z(sll_386_ML_int_3__48_) );
  MUX2_X2 sll_386_M1_2_49 ( .A(sll_386_ML_int_2__49_), .B(
        sll_386_ML_int_2__45_), .S(sll_386_n7), .Z(sll_386_ML_int_3__49_) );
  MUX2_X2 sll_386_M1_2_50 ( .A(sll_386_ML_int_2__50_), .B(
        sll_386_ML_int_2__46_), .S(sll_386_n7), .Z(sll_386_ML_int_3__50_) );
  MUX2_X2 sll_386_M1_2_51 ( .A(sll_386_ML_int_2__51_), .B(
        sll_386_ML_int_2__47_), .S(sll_386_n7), .Z(sll_386_ML_int_3__51_) );
  MUX2_X2 sll_386_M1_2_52 ( .A(sll_386_ML_int_2__52_), .B(
        sll_386_ML_int_2__48_), .S(sll_386_n7), .Z(sll_386_ML_int_3__52_) );
  MUX2_X2 sll_386_M1_3_8 ( .A(sll_386_ML_int_3__8_), .B(sll_386_ML_int_3__0_), 
        .S(div_opa_ldz_d[3]), .Z(sll_386_ML_int_4__8_) );
  MUX2_X2 sll_386_M1_3_9 ( .A(sll_386_ML_int_3__9_), .B(sll_386_ML_int_3__1_), 
        .S(div_opa_ldz_d[3]), .Z(sll_386_ML_int_4__9_) );
  MUX2_X2 sll_386_M1_3_10 ( .A(sll_386_ML_int_3__10_), .B(sll_386_ML_int_3__2_), .S(div_opa_ldz_d[3]), .Z(sll_386_ML_int_4__10_) );
  MUX2_X2 sll_386_M1_3_11 ( .A(sll_386_ML_int_3__11_), .B(sll_386_ML_int_3__3_), .S(div_opa_ldz_d[3]), .Z(sll_386_ML_int_4__11_) );
  MUX2_X2 sll_386_M1_3_12 ( .A(sll_386_ML_int_3__12_), .B(sll_386_ML_int_3__4_), .S(div_opa_ldz_d[3]), .Z(sll_386_ML_int_4__12_) );
  MUX2_X2 sll_386_M1_3_13 ( .A(sll_386_ML_int_3__13_), .B(sll_386_ML_int_3__5_), .S(div_opa_ldz_d[3]), .Z(sll_386_ML_int_4__13_) );
  MUX2_X2 sll_386_M1_3_14 ( .A(sll_386_ML_int_3__14_), .B(sll_386_ML_int_3__6_), .S(div_opa_ldz_d[3]), .Z(sll_386_ML_int_4__14_) );
  MUX2_X2 sll_386_M1_3_15 ( .A(sll_386_ML_int_3__15_), .B(sll_386_ML_int_3__7_), .S(div_opa_ldz_d[3]), .Z(sll_386_ML_int_4__15_) );
  MUX2_X2 sll_386_M1_3_16 ( .A(sll_386_ML_int_3__16_), .B(sll_386_ML_int_3__8_), .S(div_opa_ldz_d[3]), .Z(sll_386_ML_int_4__16_) );
  MUX2_X2 sll_386_M1_3_17 ( .A(sll_386_ML_int_3__17_), .B(sll_386_ML_int_3__9_), .S(div_opa_ldz_d[3]), .Z(sll_386_ML_int_4__17_) );
  MUX2_X2 sll_386_M1_3_18 ( .A(sll_386_ML_int_3__18_), .B(
        sll_386_ML_int_3__10_), .S(sll_386_n9), .Z(sll_386_ML_int_4__18_) );
  MUX2_X2 sll_386_M1_3_19 ( .A(sll_386_ML_int_3__19_), .B(
        sll_386_ML_int_3__11_), .S(div_opa_ldz_d[3]), .Z(sll_386_ML_int_4__19_) );
  MUX2_X2 sll_386_M1_3_20 ( .A(sll_386_ML_int_3__20_), .B(
        sll_386_ML_int_3__12_), .S(div_opa_ldz_d[3]), .Z(sll_386_ML_int_4__20_) );
  MUX2_X2 sll_386_M1_3_21 ( .A(sll_386_ML_int_3__21_), .B(
        sll_386_ML_int_3__13_), .S(div_opa_ldz_d[3]), .Z(sll_386_ML_int_4__21_) );
  MUX2_X2 sll_386_M1_3_22 ( .A(sll_386_ML_int_3__22_), .B(
        sll_386_ML_int_3__14_), .S(div_opa_ldz_d[3]), .Z(sll_386_ML_int_4__22_) );
  MUX2_X2 sll_386_M1_3_23 ( .A(sll_386_ML_int_3__23_), .B(
        sll_386_ML_int_3__15_), .S(div_opa_ldz_d[3]), .Z(sll_386_ML_int_4__23_) );
  MUX2_X2 sll_386_M1_3_24 ( .A(sll_386_ML_int_3__24_), .B(
        sll_386_ML_int_3__16_), .S(div_opa_ldz_d[3]), .Z(sll_386_ML_int_4__24_) );
  MUX2_X2 sll_386_M1_3_25 ( .A(sll_386_ML_int_3__25_), .B(
        sll_386_ML_int_3__17_), .S(div_opa_ldz_d[3]), .Z(sll_386_ML_int_4__25_) );
  MUX2_X2 sll_386_M1_3_26 ( .A(sll_386_ML_int_3__26_), .B(
        sll_386_ML_int_3__18_), .S(div_opa_ldz_d[3]), .Z(sll_386_ML_int_4__26_) );
  MUX2_X2 sll_386_M1_3_27 ( .A(sll_386_ML_int_3__27_), .B(
        sll_386_ML_int_3__19_), .S(div_opa_ldz_d[3]), .Z(sll_386_ML_int_4__27_) );
  MUX2_X2 sll_386_M1_3_28 ( .A(sll_386_ML_int_3__28_), .B(
        sll_386_ML_int_3__20_), .S(div_opa_ldz_d[3]), .Z(sll_386_ML_int_4__28_) );
  MUX2_X2 sll_386_M1_3_29 ( .A(sll_386_ML_int_3__29_), .B(
        sll_386_ML_int_3__21_), .S(div_opa_ldz_d[3]), .Z(sll_386_ML_int_4__29_) );
  MUX2_X2 sll_386_M1_3_30 ( .A(sll_386_ML_int_3__30_), .B(
        sll_386_ML_int_3__22_), .S(sll_386_n9), .Z(sll_386_ML_int_4__30_) );
  MUX2_X2 sll_386_M1_3_31 ( .A(sll_386_ML_int_3__31_), .B(
        sll_386_ML_int_3__23_), .S(sll_386_n9), .Z(sll_386_ML_int_4__31_) );
  MUX2_X2 sll_386_M1_3_32 ( .A(sll_386_ML_int_3__32_), .B(
        sll_386_ML_int_3__24_), .S(sll_386_n9), .Z(sll_386_ML_int_4__32_) );
  MUX2_X2 sll_386_M1_3_33 ( .A(sll_386_ML_int_3__33_), .B(
        sll_386_ML_int_3__25_), .S(sll_386_n9), .Z(sll_386_ML_int_4__33_) );
  MUX2_X2 sll_386_M1_3_34 ( .A(sll_386_ML_int_3__34_), .B(
        sll_386_ML_int_3__26_), .S(sll_386_n9), .Z(sll_386_ML_int_4__34_) );
  MUX2_X2 sll_386_M1_3_35 ( .A(sll_386_ML_int_3__35_), .B(
        sll_386_ML_int_3__27_), .S(sll_386_n9), .Z(sll_386_ML_int_4__35_) );
  MUX2_X2 sll_386_M1_3_36 ( .A(sll_386_ML_int_3__36_), .B(
        sll_386_ML_int_3__28_), .S(sll_386_n9), .Z(sll_386_ML_int_4__36_) );
  MUX2_X2 sll_386_M1_3_37 ( .A(sll_386_ML_int_3__37_), .B(
        sll_386_ML_int_3__29_), .S(sll_386_n9), .Z(sll_386_ML_int_4__37_) );
  MUX2_X2 sll_386_M1_3_38 ( .A(sll_386_ML_int_3__38_), .B(
        sll_386_ML_int_3__30_), .S(sll_386_n9), .Z(sll_386_ML_int_4__38_) );
  MUX2_X2 sll_386_M1_3_39 ( .A(sll_386_ML_int_3__39_), .B(
        sll_386_ML_int_3__31_), .S(sll_386_n9), .Z(sll_386_ML_int_4__39_) );
  MUX2_X2 sll_386_M1_3_40 ( .A(sll_386_ML_int_3__40_), .B(
        sll_386_ML_int_3__32_), .S(sll_386_n9), .Z(sll_386_ML_int_4__40_) );
  MUX2_X2 sll_386_M1_3_41 ( .A(sll_386_ML_int_3__41_), .B(
        sll_386_ML_int_3__33_), .S(sll_386_n9), .Z(sll_386_ML_int_4__41_) );
  MUX2_X2 sll_386_M1_3_42 ( .A(sll_386_ML_int_3__42_), .B(
        sll_386_ML_int_3__34_), .S(sll_386_n9), .Z(sll_386_ML_int_4__42_) );
  MUX2_X2 sll_386_M1_3_43 ( .A(sll_386_ML_int_3__43_), .B(
        sll_386_ML_int_3__35_), .S(sll_386_n9), .Z(sll_386_ML_int_4__43_) );
  MUX2_X2 sll_386_M1_3_44 ( .A(sll_386_ML_int_3__44_), .B(
        sll_386_ML_int_3__36_), .S(sll_386_n9), .Z(sll_386_ML_int_4__44_) );
  MUX2_X2 sll_386_M1_3_45 ( .A(sll_386_ML_int_3__45_), .B(
        sll_386_ML_int_3__37_), .S(sll_386_n9), .Z(sll_386_ML_int_4__45_) );
  MUX2_X2 sll_386_M1_3_46 ( .A(sll_386_ML_int_3__46_), .B(
        sll_386_ML_int_3__38_), .S(sll_386_n9), .Z(sll_386_ML_int_4__46_) );
  MUX2_X2 sll_386_M1_3_47 ( .A(sll_386_ML_int_3__47_), .B(
        sll_386_ML_int_3__39_), .S(sll_386_n9), .Z(sll_386_ML_int_4__47_) );
  MUX2_X2 sll_386_M1_3_48 ( .A(sll_386_ML_int_3__48_), .B(
        sll_386_ML_int_3__40_), .S(sll_386_n9), .Z(sll_386_ML_int_4__48_) );
  MUX2_X2 sll_386_M1_3_49 ( .A(sll_386_ML_int_3__49_), .B(
        sll_386_ML_int_3__41_), .S(sll_386_n9), .Z(sll_386_ML_int_4__49_) );
  MUX2_X2 sll_386_M1_3_50 ( .A(sll_386_ML_int_3__50_), .B(
        sll_386_ML_int_3__42_), .S(sll_386_n9), .Z(sll_386_ML_int_4__50_) );
  MUX2_X2 sll_386_M1_3_51 ( .A(sll_386_ML_int_3__51_), .B(
        sll_386_ML_int_3__43_), .S(sll_386_n9), .Z(sll_386_ML_int_4__51_) );
  MUX2_X2 sll_386_M1_3_52 ( .A(sll_386_ML_int_3__52_), .B(
        sll_386_ML_int_3__44_), .S(sll_386_n9), .Z(sll_386_ML_int_4__52_) );
  MUX2_X2 sll_386_M1_4_16 ( .A(sll_386_ML_int_4__16_), .B(sll_386_n18), .S(
        sll_386_n11), .Z(N272) );
  MUX2_X2 sll_386_M1_4_17 ( .A(sll_386_ML_int_4__17_), .B(sll_386_n17), .S(
        sll_386_n14), .Z(N273) );
  MUX2_X2 sll_386_M1_4_18 ( .A(sll_386_ML_int_4__18_), .B(sll_386_n16), .S(
        sll_386_n13), .Z(N274) );
  MUX2_X2 sll_386_M1_4_19 ( .A(sll_386_ML_int_4__19_), .B(sll_386_n15), .S(
        sll_386_n11), .Z(N275) );
  MUX2_X2 sll_386_M1_4_20 ( .A(sll_386_ML_int_4__20_), .B(sll_386_n19), .S(
        sll_386_n14), .Z(N276) );
  MUX2_X2 sll_386_M1_4_21 ( .A(sll_386_ML_int_4__21_), .B(sll_386_n20), .S(
        sll_386_n14), .Z(N277) );
  MUX2_X2 sll_386_M1_4_22 ( .A(sll_386_ML_int_4__22_), .B(sll_386_n21), .S(
        sll_386_n14), .Z(N278) );
  MUX2_X2 sll_386_M1_4_23 ( .A(sll_386_ML_int_4__23_), .B(sll_386_n22), .S(
        sll_386_n14), .Z(N279) );
  MUX2_X2 sll_386_M1_4_24 ( .A(sll_386_ML_int_4__24_), .B(sll_386_ML_int_4__8_), .S(sll_386_n14), .Z(N280) );
  MUX2_X2 sll_386_M1_4_25 ( .A(sll_386_ML_int_4__25_), .B(sll_386_ML_int_4__9_), .S(sll_386_n14), .Z(N281) );
  MUX2_X2 sll_386_M1_4_26 ( .A(sll_386_ML_int_4__26_), .B(
        sll_386_ML_int_4__10_), .S(sll_386_n14), .Z(N282) );
  MUX2_X2 sll_386_M1_4_27 ( .A(sll_386_ML_int_4__27_), .B(
        sll_386_ML_int_4__11_), .S(sll_386_n14), .Z(N283) );
  MUX2_X2 sll_386_M1_4_28 ( .A(sll_386_ML_int_4__28_), .B(
        sll_386_ML_int_4__12_), .S(sll_386_n14), .Z(N284) );
  MUX2_X2 sll_386_M1_4_29 ( .A(sll_386_ML_int_4__29_), .B(
        sll_386_ML_int_4__13_), .S(sll_386_n14), .Z(N285) );
  MUX2_X2 sll_386_M1_4_30 ( .A(sll_386_ML_int_4__30_), .B(
        sll_386_ML_int_4__14_), .S(sll_386_n14), .Z(N286) );
  MUX2_X2 sll_386_M1_4_31 ( .A(sll_386_ML_int_4__31_), .B(
        sll_386_ML_int_4__15_), .S(sll_386_n13), .Z(N287) );
  MUX2_X2 sll_386_M1_4_32 ( .A(sll_386_ML_int_4__32_), .B(
        sll_386_ML_int_4__16_), .S(sll_386_n13), .Z(N288) );
  MUX2_X2 sll_386_M1_4_33 ( .A(sll_386_ML_int_4__33_), .B(
        sll_386_ML_int_4__17_), .S(sll_386_n13), .Z(N289) );
  MUX2_X2 sll_386_M1_4_34 ( .A(sll_386_ML_int_4__34_), .B(
        sll_386_ML_int_4__18_), .S(sll_386_n13), .Z(N290) );
  MUX2_X2 sll_386_M1_4_35 ( .A(sll_386_ML_int_4__35_), .B(
        sll_386_ML_int_4__19_), .S(sll_386_n13), .Z(N291) );
  MUX2_X2 sll_386_M1_4_36 ( .A(sll_386_ML_int_4__36_), .B(
        sll_386_ML_int_4__20_), .S(sll_386_n13), .Z(N292) );
  MUX2_X2 sll_386_M1_4_37 ( .A(sll_386_ML_int_4__37_), .B(
        sll_386_ML_int_4__21_), .S(sll_386_n13), .Z(N293) );
  MUX2_X2 sll_386_M1_4_38 ( .A(sll_386_ML_int_4__38_), .B(
        sll_386_ML_int_4__22_), .S(sll_386_n13), .Z(N294) );
  MUX2_X2 sll_386_M1_4_39 ( .A(sll_386_ML_int_4__39_), .B(
        sll_386_ML_int_4__23_), .S(sll_386_n13), .Z(N295) );
  MUX2_X2 sll_386_M1_4_40 ( .A(sll_386_ML_int_4__40_), .B(
        sll_386_ML_int_4__24_), .S(sll_386_n13), .Z(N296) );
  MUX2_X2 sll_386_M1_4_41 ( .A(sll_386_ML_int_4__41_), .B(
        sll_386_ML_int_4__25_), .S(sll_386_n13), .Z(N297) );
  MUX2_X2 sll_386_M1_4_42 ( .A(sll_386_ML_int_4__42_), .B(
        sll_386_ML_int_4__26_), .S(div_opa_ldz_d[4]), .Z(N298) );
  MUX2_X2 sll_386_M1_4_43 ( .A(sll_386_ML_int_4__43_), .B(
        sll_386_ML_int_4__27_), .S(div_opa_ldz_d[4]), .Z(N299) );
  MUX2_X2 sll_386_M1_4_44 ( .A(sll_386_ML_int_4__44_), .B(
        sll_386_ML_int_4__28_), .S(div_opa_ldz_d[4]), .Z(N300) );
  MUX2_X2 sll_386_M1_4_45 ( .A(sll_386_ML_int_4__45_), .B(
        sll_386_ML_int_4__29_), .S(div_opa_ldz_d[4]), .Z(N301) );
  MUX2_X2 sll_386_M1_4_46 ( .A(sll_386_ML_int_4__46_), .B(
        sll_386_ML_int_4__30_), .S(div_opa_ldz_d[4]), .Z(N302) );
  MUX2_X2 sll_386_M1_4_47 ( .A(sll_386_ML_int_4__47_), .B(
        sll_386_ML_int_4__31_), .S(sll_386_n11), .Z(N303) );
  MUX2_X2 sll_386_M1_4_48 ( .A(sll_386_ML_int_4__48_), .B(
        sll_386_ML_int_4__32_), .S(div_opa_ldz_d[4]), .Z(N304) );
  MUX2_X2 sll_386_M1_4_49 ( .A(sll_386_ML_int_4__49_), .B(
        sll_386_ML_int_4__33_), .S(div_opa_ldz_d[4]), .Z(N305) );
  MUX2_X2 sll_386_M1_4_50 ( .A(sll_386_ML_int_4__50_), .B(
        sll_386_ML_int_4__34_), .S(div_opa_ldz_d[4]), .Z(N306) );
  MUX2_X2 sll_386_M1_4_51 ( .A(sll_386_ML_int_4__51_), .B(
        sll_386_ML_int_4__35_), .S(div_opa_ldz_d[4]), .Z(N307) );
  MUX2_X2 sll_386_M1_4_52 ( .A(sll_386_ML_int_4__52_), .B(
        sll_386_ML_int_4__36_), .S(sll_386_n11), .Z(N308) );
  NAND2_X1 r471_U180 ( .A1(fracta_mul[49]), .A2(r471_n7), .ZN(r471_n168) );
  OR2_X1 r471_U179 ( .A1(r471_n1), .A2(u6_N50), .ZN(r471_n167) );
  AND2_X1 r471_U178 ( .A1(fracta_mul[0]), .A2(r471_n56), .ZN(r471_n178) );
  OAI22_X1 r471_U177 ( .A1(fracta_mul[1]), .A2(r471_n178), .B1(r471_n178), 
        .B2(r471_n55), .ZN(r471_n177) );
  AND3_X1 r471_U176 ( .A1(r471_n168), .A2(r471_n167), .A3(r471_n177), .ZN(
        r471_n176) );
  NAND2_X1 r471_U175 ( .A1(fracta_mul[48]), .A2(r471_n8), .ZN(r471_n93) );
  NAND2_X1 r471_U174 ( .A1(fracta_mul[46]), .A2(r471_n10), .ZN(r471_n97) );
  NAND2_X1 r471_U173 ( .A1(fracta_mul[47]), .A2(r471_n9), .ZN(r471_n94) );
  AND4_X1 r471_U172 ( .A1(r471_n176), .A2(r471_n93), .A3(r471_n97), .A4(
        r471_n94), .ZN(r471_n169) );
  NAND2_X1 r471_U171 ( .A1(fracta_mul[42]), .A2(r471_n14), .ZN(r471_n105) );
  NAND2_X1 r471_U170 ( .A1(fracta_mul[41]), .A2(r471_n15), .ZN(r471_n106) );
  NAND2_X1 r471_U169 ( .A1(fracta_mul[40]), .A2(r471_n16), .ZN(r471_n109) );
  NAND2_X1 r471_U168 ( .A1(fracta_mul[39]), .A2(r471_n17), .ZN(r471_n110) );
  AND4_X1 r471_U167 ( .A1(r471_n105), .A2(r471_n106), .A3(r471_n109), .A4(
        r471_n110), .ZN(r471_n175) );
  NAND2_X1 r471_U166 ( .A1(fracta_mul[45]), .A2(r471_n11), .ZN(r471_n98) );
  NAND2_X1 r471_U165 ( .A1(fracta_mul[43]), .A2(r471_n13), .ZN(r471_n102) );
  NAND2_X1 r471_U164 ( .A1(fracta_mul[44]), .A2(r471_n12), .ZN(r471_n101) );
  AND4_X1 r471_U163 ( .A1(r471_n175), .A2(r471_n98), .A3(r471_n102), .A4(
        r471_n101), .ZN(r471_n170) );
  NAND2_X1 r471_U162 ( .A1(fracta_mul[34]), .A2(r471_n22), .ZN(r471_n121) );
  NAND2_X1 r471_U161 ( .A1(fracta_mul[33]), .A2(r471_n23), .ZN(r471_n122) );
  NAND2_X1 r471_U160 ( .A1(fracta_mul[35]), .A2(r471_n21), .ZN(r471_n118) );
  AND3_X1 r471_U159 ( .A1(r471_n121), .A2(r471_n122), .A3(r471_n118), .ZN(
        r471_n174) );
  NAND2_X1 r471_U158 ( .A1(fracta_mul[38]), .A2(r471_n18), .ZN(r471_n113) );
  NAND2_X1 r471_U157 ( .A1(fracta_mul[36]), .A2(r471_n20), .ZN(r471_n117) );
  NAND2_X1 r471_U156 ( .A1(fracta_mul[37]), .A2(r471_n19), .ZN(r471_n114) );
  AND4_X1 r471_U155 ( .A1(r471_n174), .A2(r471_n113), .A3(r471_n117), .A4(
        r471_n114), .ZN(r471_n171) );
  NAND2_X1 r471_U154 ( .A1(fracta_mul[29]), .A2(r471_n27), .ZN(r471_n130) );
  NAND2_X1 r471_U153 ( .A1(fracta_mul[28]), .A2(r471_n28), .ZN(r471_n133) );
  NAND2_X1 r471_U152 ( .A1(fracta_mul[27]), .A2(r471_n29), .ZN(r471_n134) );
  NAND2_X1 r471_U151 ( .A1(fracta_mul[26]), .A2(r471_n30), .ZN(r471_n137) );
  AND4_X1 r471_U150 ( .A1(r471_n130), .A2(r471_n133), .A3(r471_n134), .A4(
        r471_n137), .ZN(r471_n173) );
  NAND2_X1 r471_U149 ( .A1(fracta_mul[32]), .A2(r471_n24), .ZN(r471_n125) );
  NAND2_X1 r471_U148 ( .A1(fracta_mul[30]), .A2(r471_n26), .ZN(r471_n129) );
  NAND2_X1 r471_U147 ( .A1(fracta_mul[31]), .A2(r471_n25), .ZN(r471_n126) );
  AND4_X1 r471_U146 ( .A1(r471_n173), .A2(r471_n125), .A3(r471_n129), .A4(
        r471_n126), .ZN(r471_n172) );
  NAND4_X1 r471_U145 ( .A1(r471_n169), .A2(r471_n170), .A3(r471_n171), .A4(
        r471_n172), .ZN(r471_n57) );
  NAND2_X1 r471_U144 ( .A1(fracta_mul[6]), .A2(r471_n50), .ZN(r471_n158) );
  NAND2_X1 r471_U143 ( .A1(fracta_mul[4]), .A2(r471_n52), .ZN(r471_n162) );
  NAND2_X1 r471_U142 ( .A1(fracta_mul[5]), .A2(r471_n51), .ZN(r471_n159) );
  AND3_X1 r471_U141 ( .A1(r471_n158), .A2(r471_n162), .A3(r471_n159), .ZN(
        r471_n76) );
  AND2_X1 r471_U140 ( .A1(fracta_mul[51]), .A2(r471_n6), .ZN(r471_n86) );
  AND2_X1 r471_U139 ( .A1(r471_n167), .A2(r471_n168), .ZN(r471_n90) );
  NAND2_X1 r471_U138 ( .A1(fracta_mul[25]), .A2(r471_n31), .ZN(r471_n63) );
  NAND2_X1 r471_U137 ( .A1(fracta_mul[24]), .A2(r471_n32), .ZN(r471_n61) );
  NAND2_X1 r471_U136 ( .A1(fracta_mul[23]), .A2(r471_n33), .ZN(r471_n62) );
  NAND2_X1 r471_U135 ( .A1(fracta_mul[22]), .A2(r471_n34), .ZN(r471_n65) );
  NAND2_X1 r471_U134 ( .A1(fracta_mul[21]), .A2(r471_n35), .ZN(r471_n67) );
  NAND2_X1 r471_U133 ( .A1(fracta_mul[20]), .A2(r471_n36), .ZN(r471_n66) );
  NAND2_X1 r471_U132 ( .A1(fracta_mul[19]), .A2(r471_n37), .ZN(r471_n70) );
  NAND2_X1 r471_U131 ( .A1(fracta_mul[18]), .A2(r471_n38), .ZN(r471_n68) );
  NAND2_X1 r471_U130 ( .A1(fracta_mul[17]), .A2(r471_n39), .ZN(r471_n69) );
  NAND2_X1 r471_U129 ( .A1(fracta_mul[16]), .A2(r471_n40), .ZN(r471_n75) );
  NAND2_X1 r471_U128 ( .A1(fracta_mul[15]), .A2(r471_n41), .ZN(r471_n74) );
  NAND2_X1 r471_U127 ( .A1(fracta_mul[14]), .A2(r471_n42), .ZN(r471_n73) );
  NAND2_X1 r471_U126 ( .A1(fracta_mul[13]), .A2(r471_n43), .ZN(r471_n72) );
  NAND2_X1 r471_U125 ( .A1(fracta_mul[12]), .A2(r471_n44), .ZN(r471_n80) );
  NAND2_X1 r471_U124 ( .A1(fracta_mul[11]), .A2(r471_n45), .ZN(r471_n82) );
  NAND2_X1 r471_U123 ( .A1(fracta_mul[10]), .A2(r471_n46), .ZN(r471_n81) );
  NAND2_X1 r471_U122 ( .A1(fracta_mul[9]), .A2(r471_n47), .ZN(r471_n85) );
  NAND2_X1 r471_U121 ( .A1(fracta_mul[8]), .A2(r471_n48), .ZN(r471_n83) );
  NAND2_X1 r471_U120 ( .A1(fracta_mul[7]), .A2(r471_n49), .ZN(r471_n84) );
  NAND2_X1 r471_U119 ( .A1(fracta_mul[3]), .A2(r471_n53), .ZN(r471_n87) );
  NOR2_X1 r471_U118 ( .A1(r471_n56), .A2(fracta_mul[0]), .ZN(r471_n165) );
  OAI21_X1 r471_U117 ( .B1(fracta_mul[1]), .B2(r471_n5), .A(r471_n55), .ZN(
        r471_n166) );
  NAND2_X1 r471_U116 ( .A1(fracta_mul[2]), .A2(r471_n54), .ZN(r471_n88) );
  OAI211_X1 r471_U115 ( .C1(r471_n165), .C2(r471_n4), .A(r471_n166), .B(
        r471_n88), .ZN(r471_n164) );
  OAI221_X1 r471_U114 ( .B1(fracta_mul[2]), .B2(r471_n54), .C1(fracta_mul[3]), 
        .C2(r471_n53), .A(r471_n164), .ZN(r471_n163) );
  NAND3_X1 r471_U113 ( .A1(r471_n162), .A2(r471_n87), .A3(r471_n163), .ZN(
        r471_n161) );
  OAI221_X1 r471_U112 ( .B1(fracta_mul[4]), .B2(r471_n52), .C1(fracta_mul[5]), 
        .C2(r471_n51), .A(r471_n161), .ZN(r471_n160) );
  NAND3_X1 r471_U111 ( .A1(r471_n158), .A2(r471_n159), .A3(r471_n160), .ZN(
        r471_n157) );
  OAI221_X1 r471_U110 ( .B1(fracta_mul[6]), .B2(r471_n50), .C1(fracta_mul[7]), 
        .C2(r471_n49), .A(r471_n157), .ZN(r471_n156) );
  NAND3_X1 r471_U109 ( .A1(r471_n83), .A2(r471_n84), .A3(r471_n156), .ZN(
        r471_n155) );
  OAI221_X1 r471_U108 ( .B1(fracta_mul[8]), .B2(r471_n48), .C1(fracta_mul[9]), 
        .C2(r471_n47), .A(r471_n155), .ZN(r471_n154) );
  NAND3_X1 r471_U107 ( .A1(r471_n81), .A2(r471_n85), .A3(r471_n154), .ZN(
        r471_n153) );
  OAI221_X1 r471_U106 ( .B1(fracta_mul[10]), .B2(r471_n46), .C1(fracta_mul[11]), .C2(r471_n45), .A(r471_n153), .ZN(r471_n152) );
  NAND3_X1 r471_U105 ( .A1(r471_n80), .A2(r471_n82), .A3(r471_n152), .ZN(
        r471_n151) );
  OAI221_X1 r471_U104 ( .B1(fracta_mul[12]), .B2(r471_n44), .C1(fracta_mul[13]), .C2(r471_n43), .A(r471_n151), .ZN(r471_n150) );
  NAND3_X1 r471_U103 ( .A1(r471_n73), .A2(r471_n72), .A3(r471_n150), .ZN(
        r471_n149) );
  OAI221_X1 r471_U102 ( .B1(fracta_mul[14]), .B2(r471_n42), .C1(fracta_mul[15]), .C2(r471_n41), .A(r471_n149), .ZN(r471_n148) );
  NAND3_X1 r471_U101 ( .A1(r471_n75), .A2(r471_n74), .A3(r471_n148), .ZN(
        r471_n147) );
  OAI221_X1 r471_U100 ( .B1(fracta_mul[16]), .B2(r471_n40), .C1(fracta_mul[17]), .C2(r471_n39), .A(r471_n147), .ZN(r471_n146) );
  NAND3_X1 r471_U99 ( .A1(r471_n68), .A2(r471_n69), .A3(r471_n146), .ZN(
        r471_n145) );
  OAI221_X1 r471_U98 ( .B1(fracta_mul[18]), .B2(r471_n38), .C1(fracta_mul[19]), 
        .C2(r471_n37), .A(r471_n145), .ZN(r471_n144) );
  NAND3_X1 r471_U97 ( .A1(r471_n66), .A2(r471_n70), .A3(r471_n144), .ZN(
        r471_n143) );
  OAI221_X1 r471_U96 ( .B1(fracta_mul[20]), .B2(r471_n36), .C1(fracta_mul[21]), 
        .C2(r471_n35), .A(r471_n143), .ZN(r471_n142) );
  NAND3_X1 r471_U95 ( .A1(r471_n65), .A2(r471_n67), .A3(r471_n142), .ZN(
        r471_n141) );
  OAI221_X1 r471_U94 ( .B1(fracta_mul[22]), .B2(r471_n34), .C1(fracta_mul[23]), 
        .C2(r471_n33), .A(r471_n141), .ZN(r471_n140) );
  NAND3_X1 r471_U93 ( .A1(r471_n61), .A2(r471_n62), .A3(r471_n140), .ZN(
        r471_n139) );
  OAI221_X1 r471_U92 ( .B1(fracta_mul[24]), .B2(r471_n32), .C1(fracta_mul[25]), 
        .C2(r471_n31), .A(r471_n139), .ZN(r471_n138) );
  NAND3_X1 r471_U91 ( .A1(r471_n137), .A2(r471_n63), .A3(r471_n138), .ZN(
        r471_n136) );
  OAI221_X1 r471_U90 ( .B1(fracta_mul[26]), .B2(r471_n30), .C1(fracta_mul[27]), 
        .C2(r471_n29), .A(r471_n136), .ZN(r471_n135) );
  NAND3_X1 r471_U89 ( .A1(r471_n133), .A2(r471_n134), .A3(r471_n135), .ZN(
        r471_n132) );
  OAI221_X1 r471_U88 ( .B1(fracta_mul[28]), .B2(r471_n28), .C1(fracta_mul[29]), 
        .C2(r471_n27), .A(r471_n132), .ZN(r471_n131) );
  NAND3_X1 r471_U87 ( .A1(r471_n129), .A2(r471_n130), .A3(r471_n131), .ZN(
        r471_n128) );
  OAI221_X1 r471_U86 ( .B1(fracta_mul[30]), .B2(r471_n26), .C1(fracta_mul[31]), 
        .C2(r471_n25), .A(r471_n128), .ZN(r471_n127) );
  NAND3_X1 r471_U85 ( .A1(r471_n125), .A2(r471_n126), .A3(r471_n127), .ZN(
        r471_n124) );
  OAI221_X1 r471_U84 ( .B1(fracta_mul[32]), .B2(r471_n24), .C1(fracta_mul[33]), 
        .C2(r471_n23), .A(r471_n124), .ZN(r471_n123) );
  NAND3_X1 r471_U83 ( .A1(r471_n121), .A2(r471_n122), .A3(r471_n123), .ZN(
        r471_n120) );
  OAI221_X1 r471_U82 ( .B1(fracta_mul[34]), .B2(r471_n22), .C1(fracta_mul[35]), 
        .C2(r471_n21), .A(r471_n120), .ZN(r471_n119) );
  NAND3_X1 r471_U81 ( .A1(r471_n117), .A2(r471_n118), .A3(r471_n119), .ZN(
        r471_n116) );
  OAI221_X1 r471_U80 ( .B1(fracta_mul[36]), .B2(r471_n20), .C1(fracta_mul[37]), 
        .C2(r471_n19), .A(r471_n116), .ZN(r471_n115) );
  NAND3_X1 r471_U79 ( .A1(r471_n113), .A2(r471_n114), .A3(r471_n115), .ZN(
        r471_n112) );
  OAI221_X1 r471_U78 ( .B1(fracta_mul[38]), .B2(r471_n18), .C1(fracta_mul[39]), 
        .C2(r471_n17), .A(r471_n112), .ZN(r471_n111) );
  NAND3_X1 r471_U77 ( .A1(r471_n109), .A2(r471_n110), .A3(r471_n111), .ZN(
        r471_n108) );
  OAI221_X1 r471_U76 ( .B1(fracta_mul[40]), .B2(r471_n16), .C1(fracta_mul[41]), 
        .C2(r471_n15), .A(r471_n108), .ZN(r471_n107) );
  NAND3_X1 r471_U75 ( .A1(r471_n105), .A2(r471_n106), .A3(r471_n107), .ZN(
        r471_n104) );
  OAI221_X1 r471_U74 ( .B1(fracta_mul[42]), .B2(r471_n14), .C1(fracta_mul[43]), 
        .C2(r471_n13), .A(r471_n104), .ZN(r471_n103) );
  NAND3_X1 r471_U73 ( .A1(r471_n101), .A2(r471_n102), .A3(r471_n103), .ZN(
        r471_n100) );
  OAI221_X1 r471_U72 ( .B1(fracta_mul[44]), .B2(r471_n12), .C1(fracta_mul[45]), 
        .C2(r471_n11), .A(r471_n100), .ZN(r471_n99) );
  NAND3_X1 r471_U71 ( .A1(r471_n97), .A2(r471_n98), .A3(r471_n99), .ZN(
        r471_n96) );
  OAI221_X1 r471_U70 ( .B1(fracta_mul[46]), .B2(r471_n10), .C1(fracta_mul[47]), 
        .C2(r471_n9), .A(r471_n96), .ZN(r471_n95) );
  NAND3_X1 r471_U69 ( .A1(r471_n93), .A2(r471_n94), .A3(r471_n95), .ZN(
        r471_n92) );
  OAI221_X1 r471_U68 ( .B1(fracta_mul[48]), .B2(r471_n8), .C1(fracta_mul[49]), 
        .C2(r471_n7), .A(r471_n92), .ZN(r471_n91) );
  AOI22_X1 r471_U67 ( .A1(u6_N50), .A2(r471_n1), .B1(r471_n90), .B2(r471_n91), 
        .ZN(r471_n89) );
  OAI22_X1 r471_U66 ( .A1(fracta_mul[51]), .A2(r471_n6), .B1(r471_n86), .B2(
        r471_n89), .ZN(u1_N219) );
  NOR4_X1 r471_U65 ( .A1(u1_N219), .A2(r471_n86), .A3(r471_n3), .A4(r471_n2), 
        .ZN(r471_n77) );
  AND3_X1 r471_U64 ( .A1(r471_n83), .A2(r471_n84), .A3(r471_n85), .ZN(r471_n79) );
  AND4_X1 r471_U63 ( .A1(r471_n79), .A2(r471_n80), .A3(r471_n81), .A4(r471_n82), .ZN(r471_n78) );
  NAND3_X1 r471_U62 ( .A1(r471_n76), .A2(r471_n77), .A3(r471_n78), .ZN(
        r471_n58) );
  AND4_X1 r471_U61 ( .A1(r471_n72), .A2(r471_n73), .A3(r471_n74), .A4(r471_n75), .ZN(r471_n71) );
  NAND4_X1 r471_U60 ( .A1(r471_n68), .A2(r471_n69), .A3(r471_n70), .A4(
        r471_n71), .ZN(r471_n59) );
  AND3_X1 r471_U59 ( .A1(r471_n65), .A2(r471_n66), .A3(r471_n67), .ZN(r471_n64) );
  NAND4_X1 r471_U58 ( .A1(r471_n61), .A2(r471_n62), .A3(r471_n63), .A4(
        r471_n64), .ZN(r471_n60) );
  NOR4_X1 r471_U57 ( .A1(r471_n57), .A2(r471_n58), .A3(r471_n59), .A4(r471_n60), .ZN(u1_N220) );
  INV_X4 r471_U56 ( .A(u6_N0), .ZN(r471_n56) );
  INV_X4 r471_U55 ( .A(u6_N1), .ZN(r471_n55) );
  INV_X4 r471_U54 ( .A(u6_N2), .ZN(r471_n54) );
  INV_X4 r471_U53 ( .A(u6_N3), .ZN(r471_n53) );
  INV_X4 r471_U52 ( .A(u6_N4), .ZN(r471_n52) );
  INV_X4 r471_U51 ( .A(u6_N5), .ZN(r471_n51) );
  INV_X4 r471_U50 ( .A(u6_N6), .ZN(r471_n50) );
  INV_X4 r471_U49 ( .A(u6_N7), .ZN(r471_n49) );
  INV_X4 r471_U48 ( .A(u6_N8), .ZN(r471_n48) );
  INV_X4 r471_U47 ( .A(u6_N9), .ZN(r471_n47) );
  INV_X4 r471_U46 ( .A(u6_N10), .ZN(r471_n46) );
  INV_X4 r471_U45 ( .A(u6_N11), .ZN(r471_n45) );
  INV_X4 r471_U44 ( .A(u6_N12), .ZN(r471_n44) );
  INV_X4 r471_U43 ( .A(u6_N13), .ZN(r471_n43) );
  INV_X4 r471_U42 ( .A(u6_N14), .ZN(r471_n42) );
  INV_X4 r471_U41 ( .A(u6_N15), .ZN(r471_n41) );
  INV_X4 r471_U40 ( .A(u6_N16), .ZN(r471_n40) );
  INV_X4 r471_U39 ( .A(u6_N17), .ZN(r471_n39) );
  INV_X4 r471_U38 ( .A(u6_N18), .ZN(r471_n38) );
  INV_X4 r471_U37 ( .A(u6_N19), .ZN(r471_n37) );
  INV_X4 r471_U36 ( .A(u6_N20), .ZN(r471_n36) );
  INV_X4 r471_U35 ( .A(u6_N21), .ZN(r471_n35) );
  INV_X4 r471_U34 ( .A(u6_N22), .ZN(r471_n34) );
  INV_X4 r471_U33 ( .A(u6_N23), .ZN(r471_n33) );
  INV_X4 r471_U32 ( .A(u6_N24), .ZN(r471_n32) );
  INV_X4 r471_U31 ( .A(u6_N25), .ZN(r471_n31) );
  INV_X4 r471_U30 ( .A(u6_N26), .ZN(r471_n30) );
  INV_X4 r471_U29 ( .A(u6_N27), .ZN(r471_n29) );
  INV_X4 r471_U28 ( .A(u6_N28), .ZN(r471_n28) );
  INV_X4 r471_U27 ( .A(u6_N29), .ZN(r471_n27) );
  INV_X4 r471_U26 ( .A(u6_N30), .ZN(r471_n26) );
  INV_X4 r471_U25 ( .A(u6_N31), .ZN(r471_n25) );
  INV_X4 r471_U24 ( .A(u6_N32), .ZN(r471_n24) );
  INV_X4 r471_U23 ( .A(u6_N33), .ZN(r471_n23) );
  INV_X4 r471_U22 ( .A(u6_N34), .ZN(r471_n22) );
  INV_X4 r471_U21 ( .A(u6_N35), .ZN(r471_n21) );
  INV_X4 r471_U20 ( .A(u6_N36), .ZN(r471_n20) );
  INV_X4 r471_U19 ( .A(u6_N37), .ZN(r471_n19) );
  INV_X4 r471_U18 ( .A(u6_N38), .ZN(r471_n18) );
  INV_X4 r471_U17 ( .A(u6_N39), .ZN(r471_n17) );
  INV_X4 r471_U16 ( .A(u6_N40), .ZN(r471_n16) );
  INV_X4 r471_U15 ( .A(u6_N41), .ZN(r471_n15) );
  INV_X4 r471_U14 ( .A(u6_N42), .ZN(r471_n14) );
  INV_X4 r471_U13 ( .A(u6_N43), .ZN(r471_n13) );
  INV_X4 r471_U12 ( .A(u6_N44), .ZN(r471_n12) );
  INV_X4 r471_U11 ( .A(u6_N45), .ZN(r471_n11) );
  INV_X4 r471_U10 ( .A(u6_N46), .ZN(r471_n10) );
  INV_X4 r471_U9 ( .A(u6_N47), .ZN(r471_n9) );
  INV_X4 r471_U8 ( .A(u6_N48), .ZN(r471_n8) );
  INV_X4 r471_U7 ( .A(u6_N49), .ZN(r471_n7) );
  INV_X4 r471_U6 ( .A(u6_N51), .ZN(r471_n6) );
  INV_X4 r471_U5 ( .A(r471_n165), .ZN(r471_n5) );
  INV_X4 r471_U4 ( .A(fracta_mul[1]), .ZN(r471_n4) );
  INV_X4 r471_U3 ( .A(r471_n88), .ZN(r471_n3) );
  INV_X4 r471_U2 ( .A(r471_n87), .ZN(r471_n2) );
  INV_X4 r471_U1 ( .A(fracta_mul[50]), .ZN(r471_n1) );
  XOR2_X2 add_0_root_sub_0_root_u4_add_497_U7 ( .A(u4_fi_ldz_2a_0_), .B(
        u4_ldz_dif_0_), .Z(u4_div_exp3[0]) );
  XOR2_X2 add_0_root_sub_0_root_u4_add_497_U6 ( .A(u4_ldz_dif_10_), .B(
        add_0_root_sub_0_root_u4_add_497_n4), .Z(u4_div_exp3[10]) );
  XOR2_X2 add_0_root_sub_0_root_u4_add_497_U5 ( .A(u4_ldz_dif_9_), .B(
        add_0_root_sub_0_root_u4_add_497_n3), .Z(u4_div_exp3[9]) );
  AND2_X4 add_0_root_sub_0_root_u4_add_497_U4 ( .A1(u4_ldz_dif_9_), .A2(
        add_0_root_sub_0_root_u4_add_497_n3), .ZN(
        add_0_root_sub_0_root_u4_add_497_n4) );
  AND2_X4 add_0_root_sub_0_root_u4_add_497_U3 ( .A1(u4_ldz_dif_8_), .A2(
        add_0_root_sub_0_root_u4_add_497_carry_8_), .ZN(
        add_0_root_sub_0_root_u4_add_497_n3) );
  AND2_X4 add_0_root_sub_0_root_u4_add_497_U2 ( .A1(u4_fi_ldz_2a_0_), .A2(
        u4_ldz_dif_0_), .ZN(add_0_root_sub_0_root_u4_add_497_n2) );
  XOR2_X2 add_0_root_sub_0_root_u4_add_497_U1 ( .A(u4_ldz_dif_8_), .B(
        add_0_root_sub_0_root_u4_add_497_carry_8_), .Z(u4_div_exp3[8]) );
  FA_X1 add_0_root_sub_0_root_u4_add_497_U1_1 ( .A(u4_ldz_dif_1_), .B(
        u4_fi_ldz_2a_1_), .CI(add_0_root_sub_0_root_u4_add_497_n2), .CO(
        add_0_root_sub_0_root_u4_add_497_carry_2_), .S(u4_div_exp3[1]) );
  FA_X1 add_0_root_sub_0_root_u4_add_497_U1_2 ( .A(u4_ldz_dif_2_), .B(
        u4_fi_ldz_2a_2_), .CI(add_0_root_sub_0_root_u4_add_497_carry_2_), .CO(
        add_0_root_sub_0_root_u4_add_497_carry_3_), .S(u4_div_exp3[2]) );
  FA_X1 add_0_root_sub_0_root_u4_add_497_U1_3 ( .A(u4_ldz_dif_3_), .B(
        u4_fi_ldz_2a_3_), .CI(add_0_root_sub_0_root_u4_add_497_carry_3_), .CO(
        add_0_root_sub_0_root_u4_add_497_carry_4_), .S(u4_div_exp3[3]) );
  FA_X1 add_0_root_sub_0_root_u4_add_497_U1_4 ( .A(u4_ldz_dif_4_), .B(
        u4_fi_ldz_2a_4_), .CI(add_0_root_sub_0_root_u4_add_497_carry_4_), .CO(
        add_0_root_sub_0_root_u4_add_497_carry_5_), .S(u4_div_exp3[4]) );
  FA_X1 add_0_root_sub_0_root_u4_add_497_U1_5 ( .A(u4_ldz_dif_5_), .B(
        u4_fi_ldz_2a_5_), .CI(add_0_root_sub_0_root_u4_add_497_carry_5_), .CO(
        add_0_root_sub_0_root_u4_add_497_carry_6_), .S(u4_div_exp3[5]) );
  FA_X1 add_0_root_sub_0_root_u4_add_497_U1_6 ( .A(u4_ldz_dif_6_), .B(
        u4_fi_ldz_2a_6_), .CI(add_0_root_sub_0_root_u4_add_497_carry_6_), .CO(
        add_0_root_sub_0_root_u4_add_497_carry_7_), .S(u4_div_exp3[6]) );
  FA_X1 add_0_root_sub_0_root_u4_add_497_U1_7 ( .A(u4_ldz_dif_7_), .B(
        u4_fi_ldz_2a_6_), .CI(add_0_root_sub_0_root_u4_add_497_carry_7_), .CO(
        add_0_root_sub_0_root_u4_add_497_carry_8_), .S(u4_div_exp3[7]) );
  NOR2_X1 u5_mult_82_U3289 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n333), .ZN(
        u5_N0) );
  NOR2_X1 u5_mult_82_U3288 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n335), .ZN(
        u5_mult_82_ab_0__10_) );
  NOR2_X1 u5_mult_82_U3287 ( .A1(u5_mult_82_n426), .A2(u5_mult_82_n333), .ZN(
        u5_mult_82_ab_0__11_) );
  NOR2_X1 u5_mult_82_U3286 ( .A1(u5_mult_82_n424), .A2(u5_mult_82_n334), .ZN(
        u5_mult_82_ab_0__12_) );
  NOR2_X1 u5_mult_82_U3285 ( .A1(u5_mult_82_n421), .A2(u5_mult_82_n335), .ZN(
        u5_mult_82_ab_0__13_) );
  NOR2_X1 u5_mult_82_U3284 ( .A1(u5_mult_82_n418), .A2(u5_mult_82_n333), .ZN(
        u5_mult_82_ab_0__14_) );
  NOR2_X1 u5_mult_82_U3283 ( .A1(u5_mult_82_n415), .A2(u5_mult_82_n335), .ZN(
        u5_mult_82_ab_0__15_) );
  NOR2_X1 u5_mult_82_U3282 ( .A1(u5_mult_82_n412), .A2(u5_mult_82_n335), .ZN(
        u5_mult_82_ab_0__16_) );
  NOR2_X1 u5_mult_82_U3281 ( .A1(u5_mult_82_n409), .A2(u5_mult_82_n333), .ZN(
        u5_mult_82_ab_0__17_) );
  NOR2_X1 u5_mult_82_U3280 ( .A1(u5_mult_82_n476), .A2(u5_mult_82_n335), .ZN(
        u5_mult_82_ab_0__18_) );
  NOR2_X1 u5_mult_82_U3279 ( .A1(u5_mult_82_n404), .A2(u5_mult_82_n333), .ZN(
        u5_mult_82_ab_0__19_) );
  NOR2_X1 u5_mult_82_U3278 ( .A1(u5_mult_82_n443), .A2(u5_mult_82_n334), .ZN(
        u5_mult_82_ab_0__1_) );
  NOR2_X1 u5_mult_82_U3277 ( .A1(u5_mult_82_n475), .A2(u5_mult_82_n335), .ZN(
        u5_mult_82_ab_0__20_) );
  NOR2_X1 u5_mult_82_U3276 ( .A1(u5_mult_82_n402), .A2(u5_mult_82_n333), .ZN(
        u5_mult_82_ab_0__21_) );
  NOR2_X1 u5_mult_82_U3275 ( .A1(u5_mult_82_n400), .A2(u5_mult_82_n335), .ZN(
        u5_mult_82_ab_0__22_) );
  NOR2_X1 u5_mult_82_U3274 ( .A1(u5_mult_82_n398), .A2(u5_mult_82_n335), .ZN(
        u5_mult_82_ab_0__23_) );
  NOR2_X1 u5_mult_82_U3273 ( .A1(u5_mult_82_n396), .A2(u5_mult_82_n333), .ZN(
        u5_mult_82_ab_0__24_) );
  NOR2_X1 u5_mult_82_U3272 ( .A1(u5_mult_82_n394), .A2(u5_mult_82_n335), .ZN(
        u5_mult_82_ab_0__25_) );
  NOR2_X1 u5_mult_82_U3271 ( .A1(u5_mult_82_n392), .A2(u5_mult_82_n333), .ZN(
        u5_mult_82_ab_0__26_) );
  NOR2_X1 u5_mult_82_U3270 ( .A1(u5_mult_82_n390), .A2(u5_mult_82_n335), .ZN(
        u5_mult_82_ab_0__27_) );
  NOR2_X1 u5_mult_82_U3269 ( .A1(u5_mult_82_n387), .A2(u5_mult_82_n335), .ZN(
        u5_mult_82_ab_0__28_) );
  NOR2_X1 u5_mult_82_U3268 ( .A1(u5_mult_82_n386), .A2(u5_mult_82_n335), .ZN(
        u5_mult_82_ab_0__29_) );
  NOR2_X1 u5_mult_82_U3267 ( .A1(u5_mult_82_n442), .A2(u5_mult_82_n333), .ZN(
        u5_mult_82_ab_0__2_) );
  NOR2_X1 u5_mult_82_U3266 ( .A1(u5_mult_82_n384), .A2(u5_mult_82_n333), .ZN(
        u5_mult_82_ab_0__30_) );
  NOR2_X1 u5_mult_82_U3265 ( .A1(u5_mult_82_n382), .A2(u5_mult_82_n333), .ZN(
        u5_mult_82_ab_0__31_) );
  NOR2_X1 u5_mult_82_U3264 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n333), .ZN(
        u5_mult_82_ab_0__32_) );
  NOR2_X1 u5_mult_82_U3263 ( .A1(u5_mult_82_n378), .A2(u5_mult_82_n333), .ZN(
        u5_mult_82_ab_0__33_) );
  NOR2_X1 u5_mult_82_U3262 ( .A1(u5_mult_82_n376), .A2(u5_mult_82_n333), .ZN(
        u5_mult_82_ab_0__34_) );
  NOR2_X1 u5_mult_82_U3261 ( .A1(u5_mult_82_n374), .A2(u5_mult_82_n333), .ZN(
        u5_mult_82_ab_0__35_) );
  NOR2_X1 u5_mult_82_U3260 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n333), .ZN(
        u5_mult_82_ab_0__36_) );
  NOR2_X1 u5_mult_82_U3259 ( .A1(u5_mult_82_n370), .A2(u5_mult_82_n333), .ZN(
        u5_mult_82_ab_0__37_) );
  NOR2_X1 u5_mult_82_U3258 ( .A1(u5_mult_82_n368), .A2(u5_mult_82_n333), .ZN(
        u5_mult_82_ab_0__38_) );
  NOR2_X1 u5_mult_82_U3257 ( .A1(u5_mult_82_n366), .A2(u5_mult_82_n333), .ZN(
        u5_mult_82_ab_0__39_) );
  NOR2_X1 u5_mult_82_U3256 ( .A1(u5_mult_82_n478), .A2(u5_mult_82_n334), .ZN(
        u5_mult_82_ab_0__3_) );
  NOR2_X1 u5_mult_82_U3255 ( .A1(u5_mult_82_n364), .A2(u5_mult_82_n334), .ZN(
        u5_mult_82_ab_0__40_) );
  NOR2_X1 u5_mult_82_U3254 ( .A1(u5_mult_82_n362), .A2(u5_mult_82_n334), .ZN(
        u5_mult_82_ab_0__41_) );
  NOR2_X1 u5_mult_82_U3253 ( .A1(u5_mult_82_n360), .A2(u5_mult_82_n334), .ZN(
        u5_mult_82_ab_0__42_) );
  NOR2_X1 u5_mult_82_U3252 ( .A1(u5_mult_82_n356), .A2(u5_mult_82_n334), .ZN(
        u5_mult_82_ab_0__43_) );
  NOR2_X1 u5_mult_82_U3251 ( .A1(u5_mult_82_n355), .A2(u5_mult_82_n334), .ZN(
        u5_mult_82_ab_0__44_) );
  NOR2_X1 u5_mult_82_U3250 ( .A1(u5_mult_82_n352), .A2(u5_mult_82_n334), .ZN(
        u5_mult_82_ab_0__45_) );
  NOR2_X1 u5_mult_82_U3249 ( .A1(u5_mult_82_n350), .A2(u5_mult_82_n334), .ZN(
        u5_mult_82_ab_0__46_) );
  NOR2_X1 u5_mult_82_U3248 ( .A1(u5_mult_82_n348), .A2(u5_mult_82_n334), .ZN(
        u5_mult_82_ab_0__47_) );
  NOR2_X1 u5_mult_82_U3247 ( .A1(u5_mult_82_n346), .A2(u5_mult_82_n334), .ZN(
        u5_mult_82_ab_0__48_) );
  NOR2_X1 u5_mult_82_U3246 ( .A1(u5_mult_82_n343), .A2(u5_mult_82_n334), .ZN(
        u5_mult_82_ab_0__49_) );
  NOR2_X1 u5_mult_82_U3245 ( .A1(u5_mult_82_n438), .A2(u5_mult_82_n335), .ZN(
        u5_mult_82_ab_0__4_) );
  NOR2_X1 u5_mult_82_U3244 ( .A1(u5_mult_82_n342), .A2(u5_mult_82_n333), .ZN(
        u5_mult_82_ab_0__50_) );
  NOR2_X1 u5_mult_82_U3243 ( .A1(u5_mult_82_n338), .A2(u5_mult_82_n334), .ZN(
        u5_mult_82_ab_0__51_) );
  NOR2_X1 u5_mult_82_U3242 ( .A1(u5_mult_82_n336), .A2(u5_mult_82_n335), .ZN(
        u5_mult_82_ab_0__52_) );
  NOR2_X1 u5_mult_82_U3241 ( .A1(u5_mult_82_n436), .A2(u5_mult_82_n333), .ZN(
        u5_mult_82_ab_0__5_) );
  NOR2_X1 u5_mult_82_U3240 ( .A1(u5_mult_82_n434), .A2(u5_mult_82_n334), .ZN(
        u5_mult_82_ab_0__6_) );
  NOR2_X1 u5_mult_82_U3239 ( .A1(u5_mult_82_n432), .A2(u5_mult_82_n335), .ZN(
        u5_mult_82_ab_0__7_) );
  NOR2_X1 u5_mult_82_U3238 ( .A1(u5_mult_82_n430), .A2(u5_mult_82_n333), .ZN(
        u5_mult_82_ab_0__8_) );
  NOR2_X1 u5_mult_82_U3237 ( .A1(u5_mult_82_n428), .A2(u5_mult_82_n334), .ZN(
        u5_mult_82_ab_0__9_) );
  NOR2_X1 u5_mult_82_U3236 ( .A1(u5_mult_82_n480), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__0_) );
  NOR2_X1 u5_mult_82_U3235 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__10_) );
  NOR2_X1 u5_mult_82_U3234 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__11_) );
  NOR2_X1 u5_mult_82_U3233 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__12_) );
  NOR2_X1 u5_mult_82_U3232 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__13_) );
  NOR2_X1 u5_mult_82_U3231 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__14_) );
  NOR2_X1 u5_mult_82_U3230 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__15_) );
  NOR2_X1 u5_mult_82_U3229 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__16_) );
  NOR2_X1 u5_mult_82_U3228 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__17_) );
  NOR2_X1 u5_mult_82_U3227 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__18_) );
  NOR2_X1 u5_mult_82_U3226 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__19_) );
  NOR2_X1 u5_mult_82_U3225 ( .A1(u5_mult_82_n443), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__1_) );
  NOR2_X1 u5_mult_82_U3224 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__20_) );
  NOR2_X1 u5_mult_82_U3223 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__21_) );
  NOR2_X1 u5_mult_82_U3222 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__22_) );
  NOR2_X1 u5_mult_82_U3221 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__23_) );
  NOR2_X1 u5_mult_82_U3220 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__24_) );
  NOR2_X1 u5_mult_82_U3219 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__25_) );
  NOR2_X1 u5_mult_82_U3218 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__26_) );
  NOR2_X1 u5_mult_82_U3217 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__27_) );
  NOR2_X1 u5_mult_82_U3216 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__28_) );
  NOR2_X1 u5_mult_82_U3215 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__29_) );
  NOR2_X1 u5_mult_82_U3214 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n471), .ZN(
        u5_mult_82_ab_10__2_) );
  NOR2_X1 u5_mult_82_U3213 ( .A1(u5_mult_82_n384), .A2(u5_mult_82_n471), .ZN(
        u5_mult_82_ab_10__30_) );
  NOR2_X1 u5_mult_82_U3212 ( .A1(u5_mult_82_n382), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__31_) );
  NOR2_X1 u5_mult_82_U3211 ( .A1(u5_mult_82_n380), .A2(u5_mult_82_n471), .ZN(
        u5_mult_82_ab_10__32_) );
  NOR2_X1 u5_mult_82_U3210 ( .A1(u5_mult_82_n378), .A2(u5_mult_82_n471), .ZN(
        u5_mult_82_ab_10__33_) );
  NOR2_X1 u5_mult_82_U3209 ( .A1(u5_mult_82_n376), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__34_) );
  NOR2_X1 u5_mult_82_U3208 ( .A1(u5_mult_82_n374), .A2(u5_mult_82_n471), .ZN(
        u5_mult_82_ab_10__35_) );
  NOR2_X1 u5_mult_82_U3207 ( .A1(u5_mult_82_n474), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__36_) );
  NOR2_X1 u5_mult_82_U3206 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__37_) );
  NOR2_X1 u5_mult_82_U3205 ( .A1(u5_mult_82_n367), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__38_) );
  NOR2_X1 u5_mult_82_U3204 ( .A1(u5_mult_82_n366), .A2(u5_mult_82_n471), .ZN(
        u5_mult_82_ab_10__39_) );
  NOR2_X1 u5_mult_82_U3203 ( .A1(u5_mult_82_n441), .A2(u5_mult_82_n471), .ZN(
        u5_mult_82_ab_10__3_) );
  NOR2_X1 u5_mult_82_U3202 ( .A1(u5_mult_82_n364), .A2(u5_mult_82_n471), .ZN(
        u5_mult_82_ab_10__40_) );
  NOR2_X1 u5_mult_82_U3201 ( .A1(u5_mult_82_n362), .A2(u5_mult_82_n471), .ZN(
        u5_mult_82_ab_10__41_) );
  NOR2_X1 u5_mult_82_U3200 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n471), .ZN(
        u5_mult_82_ab_10__42_) );
  NOR2_X1 u5_mult_82_U3199 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n471), .ZN(
        u5_mult_82_ab_10__43_) );
  NOR2_X1 u5_mult_82_U3198 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n471), .ZN(
        u5_mult_82_ab_10__44_) );
  NOR2_X1 u5_mult_82_U3197 ( .A1(u5_mult_82_n352), .A2(u5_mult_82_n471), .ZN(
        u5_mult_82_ab_10__45_) );
  NOR2_X1 u5_mult_82_U3196 ( .A1(u5_mult_82_n350), .A2(u5_mult_82_n471), .ZN(
        u5_mult_82_ab_10__46_) );
  NOR2_X1 u5_mult_82_U3195 ( .A1(u5_mult_82_n348), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__47_) );
  NOR2_X1 u5_mult_82_U3194 ( .A1(u5_mult_82_n346), .A2(u5_mult_82_n471), .ZN(
        u5_mult_82_ab_10__48_) );
  NOR2_X1 u5_mult_82_U3193 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__49_) );
  NOR2_X1 u5_mult_82_U3192 ( .A1(u5_mult_82_n438), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__4_) );
  NOR2_X1 u5_mult_82_U3191 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__50_) );
  NOR2_X1 u5_mult_82_U3190 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__51_) );
  NOR2_X1 u5_mult_82_U3189 ( .A1(u5_mult_82_n336), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__52_) );
  NOR2_X1 u5_mult_82_U3188 ( .A1(u5_mult_82_n436), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__5_) );
  NOR2_X1 u5_mult_82_U3187 ( .A1(u5_mult_82_n434), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__6_) );
  NOR2_X1 u5_mult_82_U3186 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__7_) );
  NOR2_X1 u5_mult_82_U3185 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__8_) );
  NOR2_X1 u5_mult_82_U3184 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n309), .ZN(
        u5_mult_82_ab_10__9_) );
  NOR2_X1 u5_mult_82_U3183 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__0_) );
  NOR2_X1 u5_mult_82_U3182 ( .A1(u5_mult_82_n477), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__10_) );
  NOR2_X1 u5_mult_82_U3181 ( .A1(u5_mult_82_n426), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__11_) );
  NOR2_X1 u5_mult_82_U3180 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__12_) );
  NOR2_X1 u5_mult_82_U3179 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__13_) );
  NOR2_X1 u5_mult_82_U3178 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__14_) );
  NOR2_X1 u5_mult_82_U3177 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__15_) );
  NOR2_X1 u5_mult_82_U3176 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__16_) );
  NOR2_X1 u5_mult_82_U3175 ( .A1(u5_mult_82_n409), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__17_) );
  NOR2_X1 u5_mult_82_U3174 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__18_) );
  NOR2_X1 u5_mult_82_U3173 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__19_) );
  NOR2_X1 u5_mult_82_U3172 ( .A1(u5_mult_82_n443), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__1_) );
  NOR2_X1 u5_mult_82_U3171 ( .A1(u5_mult_82_n475), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__20_) );
  NOR2_X1 u5_mult_82_U3170 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__21_) );
  NOR2_X1 u5_mult_82_U3169 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__22_) );
  NOR2_X1 u5_mult_82_U3168 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__23_) );
  NOR2_X1 u5_mult_82_U3167 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__24_) );
  NOR2_X1 u5_mult_82_U3166 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__25_) );
  NOR2_X1 u5_mult_82_U3165 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__26_) );
  NOR2_X1 u5_mult_82_U3164 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__27_) );
  NOR2_X1 u5_mult_82_U3163 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__28_) );
  NOR2_X1 u5_mult_82_U3162 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__29_) );
  NOR2_X1 u5_mult_82_U3161 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n470), .ZN(
        u5_mult_82_ab_11__2_) );
  NOR2_X1 u5_mult_82_U3160 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n470), .ZN(
        u5_mult_82_ab_11__30_) );
  NOR2_X1 u5_mult_82_U3159 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n470), .ZN(
        u5_mult_82_ab_11__31_) );
  NOR2_X1 u5_mult_82_U3158 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__32_) );
  NOR2_X1 u5_mult_82_U3157 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n470), .ZN(
        u5_mult_82_ab_11__33_) );
  NOR2_X1 u5_mult_82_U3156 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__34_) );
  NOR2_X1 u5_mult_82_U3155 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__35_) );
  NOR2_X1 u5_mult_82_U3154 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__36_) );
  NOR2_X1 u5_mult_82_U3153 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__37_) );
  NOR2_X1 u5_mult_82_U3152 ( .A1(u5_mult_82_n367), .A2(u5_mult_82_n470), .ZN(
        u5_mult_82_ab_11__38_) );
  NOR2_X1 u5_mult_82_U3151 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n470), .ZN(
        u5_mult_82_ab_11__39_) );
  NOR2_X1 u5_mult_82_U3150 ( .A1(u5_mult_82_n441), .A2(u5_mult_82_n470), .ZN(
        u5_mult_82_ab_11__3_) );
  NOR2_X1 u5_mult_82_U3149 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n470), .ZN(
        u5_mult_82_ab_11__40_) );
  NOR2_X1 u5_mult_82_U3148 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n470), .ZN(
        u5_mult_82_ab_11__41_) );
  NOR2_X1 u5_mult_82_U3147 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n470), .ZN(
        u5_mult_82_ab_11__42_) );
  NOR2_X1 u5_mult_82_U3146 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n470), .ZN(
        u5_mult_82_ab_11__43_) );
  NOR2_X1 u5_mult_82_U3145 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n470), .ZN(
        u5_mult_82_ab_11__44_) );
  NOR2_X1 u5_mult_82_U3144 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n470), .ZN(
        u5_mult_82_ab_11__45_) );
  NOR2_X1 u5_mult_82_U3143 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__46_) );
  NOR2_X1 u5_mult_82_U3142 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__47_) );
  NOR2_X1 u5_mult_82_U3141 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n470), .ZN(
        u5_mult_82_ab_11__48_) );
  NOR2_X1 u5_mult_82_U3140 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__49_) );
  NOR2_X1 u5_mult_82_U3139 ( .A1(u5_mult_82_n438), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__4_) );
  NOR2_X1 u5_mult_82_U3138 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__50_) );
  NOR2_X1 u5_mult_82_U3137 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__51_) );
  NOR2_X1 u5_mult_82_U3136 ( .A1(u5_mult_82_n336), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__52_) );
  NOR2_X1 u5_mult_82_U3135 ( .A1(u5_mult_82_n436), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__5_) );
  NOR2_X1 u5_mult_82_U3134 ( .A1(u5_mult_82_n434), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__6_) );
  NOR2_X1 u5_mult_82_U3133 ( .A1(u5_mult_82_n432), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__7_) );
  NOR2_X1 u5_mult_82_U3132 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__8_) );
  NOR2_X1 u5_mult_82_U3131 ( .A1(u5_mult_82_n428), .A2(u5_mult_82_n308), .ZN(
        u5_mult_82_ab_11__9_) );
  NOR2_X1 u5_mult_82_U3130 ( .A1(u5_mult_82_n480), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__0_) );
  NOR2_X1 u5_mult_82_U3129 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__10_) );
  NOR2_X1 u5_mult_82_U3128 ( .A1(u5_mult_82_n426), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__11_) );
  NOR2_X1 u5_mult_82_U3127 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__12_) );
  NOR2_X1 u5_mult_82_U3126 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__13_) );
  NOR2_X1 u5_mult_82_U3125 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__14_) );
  NOR2_X1 u5_mult_82_U3124 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__15_) );
  NOR2_X1 u5_mult_82_U3123 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__16_) );
  NOR2_X1 u5_mult_82_U3122 ( .A1(u5_mult_82_n409), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__17_) );
  NOR2_X1 u5_mult_82_U3121 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__18_) );
  NOR2_X1 u5_mult_82_U3120 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__19_) );
  NOR2_X1 u5_mult_82_U3119 ( .A1(u5_mult_82_n443), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__1_) );
  NOR2_X1 u5_mult_82_U3118 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__20_) );
  NOR2_X1 u5_mult_82_U3117 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__21_) );
  NOR2_X1 u5_mult_82_U3116 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__22_) );
  NOR2_X1 u5_mult_82_U3115 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__23_) );
  NOR2_X1 u5_mult_82_U3114 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__24_) );
  NOR2_X1 u5_mult_82_U3113 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__25_) );
  NOR2_X1 u5_mult_82_U3112 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__26_) );
  NOR2_X1 u5_mult_82_U3111 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__27_) );
  NOR2_X1 u5_mult_82_U3110 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__28_) );
  NOR2_X1 u5_mult_82_U3109 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__29_) );
  NOR2_X1 u5_mult_82_U3108 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__2_) );
  NOR2_X1 u5_mult_82_U3107 ( .A1(u5_mult_82_n384), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__30_) );
  NOR2_X1 u5_mult_82_U3106 ( .A1(u5_mult_82_n382), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__31_) );
  NOR2_X1 u5_mult_82_U3105 ( .A1(u5_mult_82_n380), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__32_) );
  NOR2_X1 u5_mult_82_U3104 ( .A1(u5_mult_82_n378), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__33_) );
  NOR2_X1 u5_mult_82_U3103 ( .A1(u5_mult_82_n376), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__34_) );
  NOR2_X1 u5_mult_82_U3102 ( .A1(u5_mult_82_n374), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__35_) );
  NOR2_X1 u5_mult_82_U3101 ( .A1(u5_mult_82_n474), .A2(u5_mult_82_n307), .ZN(
        u5_mult_82_ab_12__36_) );
  NOR2_X1 u5_mult_82_U3100 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n307), .ZN(
        u5_mult_82_ab_12__37_) );
  NOR2_X1 u5_mult_82_U3099 ( .A1(u5_mult_82_n367), .A2(u5_mult_82_n307), .ZN(
        u5_mult_82_ab_12__38_) );
  NOR2_X1 u5_mult_82_U3098 ( .A1(u5_mult_82_n366), .A2(u5_mult_82_n307), .ZN(
        u5_mult_82_ab_12__39_) );
  NOR2_X1 u5_mult_82_U3097 ( .A1(u5_mult_82_n441), .A2(u5_mult_82_n307), .ZN(
        u5_mult_82_ab_12__3_) );
  NOR2_X1 u5_mult_82_U3096 ( .A1(u5_mult_82_n364), .A2(u5_mult_82_n307), .ZN(
        u5_mult_82_ab_12__40_) );
  NOR2_X1 u5_mult_82_U3095 ( .A1(u5_mult_82_n362), .A2(u5_mult_82_n307), .ZN(
        u5_mult_82_ab_12__41_) );
  NOR2_X1 u5_mult_82_U3094 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n307), .ZN(
        u5_mult_82_ab_12__42_) );
  NOR2_X1 u5_mult_82_U3093 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n307), .ZN(
        u5_mult_82_ab_12__43_) );
  NOR2_X1 u5_mult_82_U3092 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n307), .ZN(
        u5_mult_82_ab_12__44_) );
  NOR2_X1 u5_mult_82_U3091 ( .A1(u5_mult_82_n352), .A2(u5_mult_82_n307), .ZN(
        u5_mult_82_ab_12__45_) );
  NOR2_X1 u5_mult_82_U3090 ( .A1(u5_mult_82_n350), .A2(u5_mult_82_n307), .ZN(
        u5_mult_82_ab_12__46_) );
  NOR2_X1 u5_mult_82_U3089 ( .A1(u5_mult_82_n348), .A2(u5_mult_82_n307), .ZN(
        u5_mult_82_ab_12__47_) );
  NOR2_X1 u5_mult_82_U3088 ( .A1(u5_mult_82_n346), .A2(u5_mult_82_n307), .ZN(
        u5_mult_82_ab_12__48_) );
  NOR2_X1 u5_mult_82_U3087 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n307), .ZN(
        u5_mult_82_ab_12__49_) );
  NOR2_X1 u5_mult_82_U3086 ( .A1(u5_mult_82_n438), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__4_) );
  NOR2_X1 u5_mult_82_U3085 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__50_) );
  NOR2_X1 u5_mult_82_U3084 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__51_) );
  NOR2_X1 u5_mult_82_U3083 ( .A1(u5_mult_82_n336), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__52_) );
  NOR2_X1 u5_mult_82_U3082 ( .A1(u5_mult_82_n436), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__5_) );
  NOR2_X1 u5_mult_82_U3081 ( .A1(u5_mult_82_n434), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__6_) );
  NOR2_X1 u5_mult_82_U3080 ( .A1(u5_mult_82_n432), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__7_) );
  NOR2_X1 u5_mult_82_U3079 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__8_) );
  NOR2_X1 u5_mult_82_U3078 ( .A1(u5_mult_82_n428), .A2(u5_mult_82_n306), .ZN(
        u5_mult_82_ab_12__9_) );
  NOR2_X1 u5_mult_82_U3077 ( .A1(u5_mult_82_n480), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__0_) );
  NOR2_X1 u5_mult_82_U3076 ( .A1(u5_mult_82_n477), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__10_) );
  NOR2_X1 u5_mult_82_U3075 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__11_) );
  NOR2_X1 u5_mult_82_U3074 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__12_) );
  NOR2_X1 u5_mult_82_U3073 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__13_) );
  NOR2_X1 u5_mult_82_U3072 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__14_) );
  NOR2_X1 u5_mult_82_U3071 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__15_) );
  NOR2_X1 u5_mult_82_U3070 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__16_) );
  NOR2_X1 u5_mult_82_U3069 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__17_) );
  NOR2_X1 u5_mult_82_U3068 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__18_) );
  NOR2_X1 u5_mult_82_U3067 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__19_) );
  NOR2_X1 u5_mult_82_U3066 ( .A1(u5_mult_82_n443), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__1_) );
  NOR2_X1 u5_mult_82_U3065 ( .A1(u5_mult_82_n475), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__20_) );
  NOR2_X1 u5_mult_82_U3064 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__21_) );
  NOR2_X1 u5_mult_82_U3063 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__22_) );
  NOR2_X1 u5_mult_82_U3062 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__23_) );
  NOR2_X1 u5_mult_82_U3061 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__24_) );
  NOR2_X1 u5_mult_82_U3060 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__25_) );
  NOR2_X1 u5_mult_82_U3059 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__26_) );
  NOR2_X1 u5_mult_82_U3058 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__27_) );
  NOR2_X1 u5_mult_82_U3057 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__28_) );
  NOR2_X1 u5_mult_82_U3056 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__29_) );
  NOR2_X1 u5_mult_82_U3055 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__2_) );
  NOR2_X1 u5_mult_82_U3054 ( .A1(u5_mult_82_n384), .A2(u5_mult_82_n305), .ZN(
        u5_mult_82_ab_13__30_) );
  NOR2_X1 u5_mult_82_U3053 ( .A1(u5_mult_82_n382), .A2(u5_mult_82_n305), .ZN(
        u5_mult_82_ab_13__31_) );
  NOR2_X1 u5_mult_82_U3052 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n305), .ZN(
        u5_mult_82_ab_13__32_) );
  NOR2_X1 u5_mult_82_U3051 ( .A1(u5_mult_82_n378), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__33_) );
  NOR2_X1 u5_mult_82_U3050 ( .A1(u5_mult_82_n376), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__34_) );
  NOR2_X1 u5_mult_82_U3049 ( .A1(u5_mult_82_n374), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__35_) );
  NOR2_X1 u5_mult_82_U3048 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n305), .ZN(
        u5_mult_82_ab_13__36_) );
  NOR2_X1 u5_mult_82_U3047 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n305), .ZN(
        u5_mult_82_ab_13__37_) );
  NOR2_X1 u5_mult_82_U3046 ( .A1(u5_mult_82_n367), .A2(u5_mult_82_n305), .ZN(
        u5_mult_82_ab_13__38_) );
  NOR2_X1 u5_mult_82_U3045 ( .A1(u5_mult_82_n366), .A2(u5_mult_82_n305), .ZN(
        u5_mult_82_ab_13__39_) );
  NOR2_X1 u5_mult_82_U3044 ( .A1(u5_mult_82_n441), .A2(u5_mult_82_n305), .ZN(
        u5_mult_82_ab_13__3_) );
  NOR2_X1 u5_mult_82_U3043 ( .A1(u5_mult_82_n364), .A2(u5_mult_82_n305), .ZN(
        u5_mult_82_ab_13__40_) );
  NOR2_X1 u5_mult_82_U3042 ( .A1(u5_mult_82_n362), .A2(u5_mult_82_n305), .ZN(
        u5_mult_82_ab_13__41_) );
  NOR2_X1 u5_mult_82_U3041 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n305), .ZN(
        u5_mult_82_ab_13__42_) );
  NOR2_X1 u5_mult_82_U3040 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n305), .ZN(
        u5_mult_82_ab_13__43_) );
  NOR2_X1 u5_mult_82_U3039 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n305), .ZN(
        u5_mult_82_ab_13__44_) );
  NOR2_X1 u5_mult_82_U3038 ( .A1(u5_mult_82_n352), .A2(u5_mult_82_n305), .ZN(
        u5_mult_82_ab_13__45_) );
  NOR2_X1 u5_mult_82_U3037 ( .A1(u5_mult_82_n350), .A2(u5_mult_82_n305), .ZN(
        u5_mult_82_ab_13__46_) );
  NOR2_X1 u5_mult_82_U3036 ( .A1(u5_mult_82_n348), .A2(u5_mult_82_n305), .ZN(
        u5_mult_82_ab_13__47_) );
  NOR2_X1 u5_mult_82_U3035 ( .A1(u5_mult_82_n346), .A2(u5_mult_82_n305), .ZN(
        u5_mult_82_ab_13__48_) );
  NOR2_X1 u5_mult_82_U3034 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n305), .ZN(
        u5_mult_82_ab_13__49_) );
  NOR2_X1 u5_mult_82_U3033 ( .A1(u5_mult_82_n438), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__4_) );
  NOR2_X1 u5_mult_82_U3032 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__50_) );
  NOR2_X1 u5_mult_82_U3031 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__51_) );
  NOR2_X1 u5_mult_82_U3030 ( .A1(u5_mult_82_n336), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__52_) );
  NOR2_X1 u5_mult_82_U3029 ( .A1(u5_mult_82_n436), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__5_) );
  NOR2_X1 u5_mult_82_U3028 ( .A1(u5_mult_82_n434), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__6_) );
  NOR2_X1 u5_mult_82_U3027 ( .A1(u5_mult_82_n432), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__7_) );
  NOR2_X1 u5_mult_82_U3026 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__8_) );
  NOR2_X1 u5_mult_82_U3025 ( .A1(u5_mult_82_n428), .A2(u5_mult_82_n304), .ZN(
        u5_mult_82_ab_13__9_) );
  NOR2_X1 u5_mult_82_U3024 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__0_) );
  NOR2_X1 u5_mult_82_U3023 ( .A1(u5_mult_82_n477), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__10_) );
  NOR2_X1 u5_mult_82_U3022 ( .A1(u5_mult_82_n426), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__11_) );
  NOR2_X1 u5_mult_82_U3021 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__12_) );
  NOR2_X1 u5_mult_82_U3020 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__13_) );
  NOR2_X1 u5_mult_82_U3019 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__14_) );
  NOR2_X1 u5_mult_82_U3018 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__15_) );
  NOR2_X1 u5_mult_82_U3017 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__16_) );
  NOR2_X1 u5_mult_82_U3016 ( .A1(u5_mult_82_n409), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__17_) );
  NOR2_X1 u5_mult_82_U3015 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__18_) );
  NOR2_X1 u5_mult_82_U3014 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__19_) );
  NOR2_X1 u5_mult_82_U3013 ( .A1(u5_mult_82_n443), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__1_) );
  NOR2_X1 u5_mult_82_U3012 ( .A1(u5_mult_82_n475), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__20_) );
  NOR2_X1 u5_mult_82_U3011 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__21_) );
  NOR2_X1 u5_mult_82_U3010 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__22_) );
  NOR2_X1 u5_mult_82_U3009 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__23_) );
  NOR2_X1 u5_mult_82_U3008 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__24_) );
  NOR2_X1 u5_mult_82_U3007 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__25_) );
  NOR2_X1 u5_mult_82_U3006 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__26_) );
  NOR2_X1 u5_mult_82_U3005 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__27_) );
  NOR2_X1 u5_mult_82_U3004 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__28_) );
  NOR2_X1 u5_mult_82_U3003 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__29_) );
  NOR2_X1 u5_mult_82_U3002 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__2_) );
  NOR2_X1 u5_mult_82_U3001 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__30_) );
  NOR2_X1 u5_mult_82_U3000 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__31_) );
  NOR2_X1 u5_mult_82_U2999 ( .A1(u5_mult_82_n380), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__32_) );
  NOR2_X1 u5_mult_82_U2998 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__33_) );
  NOR2_X1 u5_mult_82_U2997 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__34_) );
  NOR2_X1 u5_mult_82_U2996 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__35_) );
  NOR2_X1 u5_mult_82_U2995 ( .A1(u5_mult_82_n474), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__36_) );
  NOR2_X1 u5_mult_82_U2994 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__37_) );
  NOR2_X1 u5_mult_82_U2993 ( .A1(u5_mult_82_n367), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__38_) );
  NOR2_X1 u5_mult_82_U2992 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__39_) );
  NOR2_X1 u5_mult_82_U2991 ( .A1(u5_mult_82_n441), .A2(u5_mult_82_n469), .ZN(
        u5_mult_82_ab_14__3_) );
  NOR2_X1 u5_mult_82_U2990 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__40_) );
  NOR2_X1 u5_mult_82_U2989 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n469), .ZN(
        u5_mult_82_ab_14__41_) );
  NOR2_X1 u5_mult_82_U2988 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n469), .ZN(
        u5_mult_82_ab_14__42_) );
  NOR2_X1 u5_mult_82_U2987 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n469), .ZN(
        u5_mult_82_ab_14__43_) );
  NOR2_X1 u5_mult_82_U2986 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n469), .ZN(
        u5_mult_82_ab_14__44_) );
  NOR2_X1 u5_mult_82_U2985 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n469), .ZN(
        u5_mult_82_ab_14__45_) );
  NOR2_X1 u5_mult_82_U2984 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n469), .ZN(
        u5_mult_82_ab_14__46_) );
  NOR2_X1 u5_mult_82_U2983 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n469), .ZN(
        u5_mult_82_ab_14__47_) );
  NOR2_X1 u5_mult_82_U2982 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n469), .ZN(
        u5_mult_82_ab_14__48_) );
  NOR2_X1 u5_mult_82_U2981 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n469), .ZN(
        u5_mult_82_ab_14__49_) );
  NOR2_X1 u5_mult_82_U2980 ( .A1(u5_mult_82_n438), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__4_) );
  NOR2_X1 u5_mult_82_U2979 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__50_) );
  NOR2_X1 u5_mult_82_U2978 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__51_) );
  NOR2_X1 u5_mult_82_U2977 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__52_) );
  NOR2_X1 u5_mult_82_U2976 ( .A1(u5_mult_82_n436), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__5_) );
  NOR2_X1 u5_mult_82_U2975 ( .A1(u5_mult_82_n434), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__6_) );
  NOR2_X1 u5_mult_82_U2974 ( .A1(u5_mult_82_n432), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__7_) );
  NOR2_X1 u5_mult_82_U2973 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__8_) );
  NOR2_X1 u5_mult_82_U2972 ( .A1(u5_mult_82_n428), .A2(u5_mult_82_n303), .ZN(
        u5_mult_82_ab_14__9_) );
  NOR2_X1 u5_mult_82_U2971 ( .A1(u5_mult_82_n480), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__0_) );
  NOR2_X1 u5_mult_82_U2970 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__10_) );
  NOR2_X1 u5_mult_82_U2969 ( .A1(u5_mult_82_n426), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__11_) );
  NOR2_X1 u5_mult_82_U2968 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__12_) );
  NOR2_X1 u5_mult_82_U2967 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__13_) );
  NOR2_X1 u5_mult_82_U2966 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__14_) );
  NOR2_X1 u5_mult_82_U2965 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__15_) );
  NOR2_X1 u5_mult_82_U2964 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__16_) );
  NOR2_X1 u5_mult_82_U2963 ( .A1(u5_mult_82_n409), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__17_) );
  NOR2_X1 u5_mult_82_U2962 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__18_) );
  NOR2_X1 u5_mult_82_U2961 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__19_) );
  NOR2_X1 u5_mult_82_U2960 ( .A1(u5_mult_82_n443), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__1_) );
  NOR2_X1 u5_mult_82_U2959 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__20_) );
  NOR2_X1 u5_mult_82_U2958 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__21_) );
  NOR2_X1 u5_mult_82_U2957 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__22_) );
  NOR2_X1 u5_mult_82_U2956 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__23_) );
  NOR2_X1 u5_mult_82_U2955 ( .A1(u5_mult_82_n396), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__24_) );
  NOR2_X1 u5_mult_82_U2954 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__25_) );
  NOR2_X1 u5_mult_82_U2953 ( .A1(u5_mult_82_n392), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__26_) );
  NOR2_X1 u5_mult_82_U2952 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__27_) );
  NOR2_X1 u5_mult_82_U2951 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__28_) );
  NOR2_X1 u5_mult_82_U2950 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__29_) );
  NOR2_X1 u5_mult_82_U2949 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__2_) );
  NOR2_X1 u5_mult_82_U2948 ( .A1(u5_mult_82_n384), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__30_) );
  NOR2_X1 u5_mult_82_U2947 ( .A1(u5_mult_82_n382), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__31_) );
  NOR2_X1 u5_mult_82_U2946 ( .A1(u5_mult_82_n380), .A2(u5_mult_82_n468), .ZN(
        u5_mult_82_ab_15__32_) );
  NOR2_X1 u5_mult_82_U2945 ( .A1(u5_mult_82_n378), .A2(u5_mult_82_n468), .ZN(
        u5_mult_82_ab_15__33_) );
  NOR2_X1 u5_mult_82_U2944 ( .A1(u5_mult_82_n376), .A2(u5_mult_82_n468), .ZN(
        u5_mult_82_ab_15__34_) );
  NOR2_X1 u5_mult_82_U2943 ( .A1(u5_mult_82_n374), .A2(u5_mult_82_n302), .ZN(
        u5_mult_82_ab_15__35_) );
  NOR2_X1 u5_mult_82_U2942 ( .A1(u5_mult_82_n474), .A2(u5_mult_82_n302), .ZN(
        u5_mult_82_ab_15__36_) );
  NOR2_X1 u5_mult_82_U2941 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n302), .ZN(
        u5_mult_82_ab_15__37_) );
  NOR2_X1 u5_mult_82_U2940 ( .A1(u5_mult_82_n367), .A2(u5_mult_82_n302), .ZN(
        u5_mult_82_ab_15__38_) );
  NOR2_X1 u5_mult_82_U2939 ( .A1(u5_mult_82_n366), .A2(u5_mult_82_n468), .ZN(
        u5_mult_82_ab_15__39_) );
  NOR2_X1 u5_mult_82_U2938 ( .A1(u5_mult_82_n441), .A2(u5_mult_82_n302), .ZN(
        u5_mult_82_ab_15__3_) );
  NOR2_X1 u5_mult_82_U2937 ( .A1(u5_mult_82_n364), .A2(u5_mult_82_n302), .ZN(
        u5_mult_82_ab_15__40_) );
  NOR2_X1 u5_mult_82_U2936 ( .A1(u5_mult_82_n362), .A2(u5_mult_82_n302), .ZN(
        u5_mult_82_ab_15__41_) );
  NOR2_X1 u5_mult_82_U2935 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n302), .ZN(
        u5_mult_82_ab_15__42_) );
  NOR2_X1 u5_mult_82_U2934 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n302), .ZN(
        u5_mult_82_ab_15__43_) );
  NOR2_X1 u5_mult_82_U2933 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n302), .ZN(
        u5_mult_82_ab_15__44_) );
  NOR2_X1 u5_mult_82_U2932 ( .A1(u5_mult_82_n352), .A2(u5_mult_82_n302), .ZN(
        u5_mult_82_ab_15__45_) );
  NOR2_X1 u5_mult_82_U2931 ( .A1(u5_mult_82_n350), .A2(u5_mult_82_n302), .ZN(
        u5_mult_82_ab_15__46_) );
  NOR2_X1 u5_mult_82_U2930 ( .A1(u5_mult_82_n348), .A2(u5_mult_82_n302), .ZN(
        u5_mult_82_ab_15__47_) );
  NOR2_X1 u5_mult_82_U2929 ( .A1(u5_mult_82_n346), .A2(u5_mult_82_n302), .ZN(
        u5_mult_82_ab_15__48_) );
  NOR2_X1 u5_mult_82_U2928 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n302), .ZN(
        u5_mult_82_ab_15__49_) );
  NOR2_X1 u5_mult_82_U2927 ( .A1(u5_mult_82_n438), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__4_) );
  NOR2_X1 u5_mult_82_U2926 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__50_) );
  NOR2_X1 u5_mult_82_U2925 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__51_) );
  NOR2_X1 u5_mult_82_U2924 ( .A1(u5_mult_82_n336), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__52_) );
  NOR2_X1 u5_mult_82_U2923 ( .A1(u5_mult_82_n436), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__5_) );
  NOR2_X1 u5_mult_82_U2922 ( .A1(u5_mult_82_n434), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__6_) );
  NOR2_X1 u5_mult_82_U2921 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__7_) );
  NOR2_X1 u5_mult_82_U2920 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__8_) );
  NOR2_X1 u5_mult_82_U2919 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n301), .ZN(
        u5_mult_82_ab_15__9_) );
  NOR2_X1 u5_mult_82_U2918 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__0_) );
  NOR2_X1 u5_mult_82_U2917 ( .A1(u5_mult_82_n477), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__10_) );
  NOR2_X1 u5_mult_82_U2916 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__11_) );
  NOR2_X1 u5_mult_82_U2915 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__12_) );
  NOR2_X1 u5_mult_82_U2914 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__13_) );
  NOR2_X1 u5_mult_82_U2913 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__14_) );
  NOR2_X1 u5_mult_82_U2912 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__15_) );
  NOR2_X1 u5_mult_82_U2911 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__16_) );
  NOR2_X1 u5_mult_82_U2910 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__17_) );
  NOR2_X1 u5_mult_82_U2909 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__18_) );
  NOR2_X1 u5_mult_82_U2908 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__19_) );
  NOR2_X1 u5_mult_82_U2907 ( .A1(u5_mult_82_n443), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__1_) );
  NOR2_X1 u5_mult_82_U2906 ( .A1(u5_mult_82_n475), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__20_) );
  NOR2_X1 u5_mult_82_U2905 ( .A1(u5_mult_82_n402), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__21_) );
  NOR2_X1 u5_mult_82_U2904 ( .A1(u5_mult_82_n400), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__22_) );
  NOR2_X1 u5_mult_82_U2903 ( .A1(u5_mult_82_n398), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__23_) );
  NOR2_X1 u5_mult_82_U2902 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__24_) );
  NOR2_X1 u5_mult_82_U2901 ( .A1(u5_mult_82_n394), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__25_) );
  NOR2_X1 u5_mult_82_U2900 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__26_) );
  NOR2_X1 u5_mult_82_U2899 ( .A1(u5_mult_82_n390), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__27_) );
  NOR2_X1 u5_mult_82_U2898 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__28_) );
  NOR2_X1 u5_mult_82_U2897 ( .A1(u5_mult_82_n386), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__29_) );
  NOR2_X1 u5_mult_82_U2896 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n300), .ZN(
        u5_mult_82_ab_16__2_) );
  NOR2_X1 u5_mult_82_U2895 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n300), .ZN(
        u5_mult_82_ab_16__30_) );
  NOR2_X1 u5_mult_82_U2894 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n300), .ZN(
        u5_mult_82_ab_16__31_) );
  NOR2_X1 u5_mult_82_U2893 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n300), .ZN(
        u5_mult_82_ab_16__32_) );
  NOR2_X1 u5_mult_82_U2892 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n300), .ZN(
        u5_mult_82_ab_16__33_) );
  NOR2_X1 u5_mult_82_U2891 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n300), .ZN(
        u5_mult_82_ab_16__34_) );
  NOR2_X1 u5_mult_82_U2890 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n300), .ZN(
        u5_mult_82_ab_16__35_) );
  NOR2_X1 u5_mult_82_U2889 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n467), .ZN(
        u5_mult_82_ab_16__36_) );
  NOR2_X1 u5_mult_82_U2888 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n467), .ZN(
        u5_mult_82_ab_16__37_) );
  NOR2_X1 u5_mult_82_U2887 ( .A1(u5_mult_82_n367), .A2(u5_mult_82_n467), .ZN(
        u5_mult_82_ab_16__38_) );
  NOR2_X1 u5_mult_82_U2886 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n467), .ZN(
        u5_mult_82_ab_16__39_) );
  NOR2_X1 u5_mult_82_U2885 ( .A1(u5_mult_82_n441), .A2(u5_mult_82_n300), .ZN(
        u5_mult_82_ab_16__3_) );
  NOR2_X1 u5_mult_82_U2884 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n300), .ZN(
        u5_mult_82_ab_16__40_) );
  NOR2_X1 u5_mult_82_U2883 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n300), .ZN(
        u5_mult_82_ab_16__41_) );
  NOR2_X1 u5_mult_82_U2882 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n300), .ZN(
        u5_mult_82_ab_16__42_) );
  NOR2_X1 u5_mult_82_U2881 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n300), .ZN(
        u5_mult_82_ab_16__43_) );
  NOR2_X1 u5_mult_82_U2880 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n300), .ZN(
        u5_mult_82_ab_16__44_) );
  NOR2_X1 u5_mult_82_U2879 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n300), .ZN(
        u5_mult_82_ab_16__45_) );
  NOR2_X1 u5_mult_82_U2878 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n300), .ZN(
        u5_mult_82_ab_16__46_) );
  NOR2_X1 u5_mult_82_U2877 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n300), .ZN(
        u5_mult_82_ab_16__47_) );
  NOR2_X1 u5_mult_82_U2876 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n300), .ZN(
        u5_mult_82_ab_16__48_) );
  NOR2_X1 u5_mult_82_U2875 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n300), .ZN(
        u5_mult_82_ab_16__49_) );
  NOR2_X1 u5_mult_82_U2874 ( .A1(u5_mult_82_n438), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__4_) );
  NOR2_X1 u5_mult_82_U2873 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__50_) );
  NOR2_X1 u5_mult_82_U2872 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__51_) );
  NOR2_X1 u5_mult_82_U2871 ( .A1(u5_mult_82_n336), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__52_) );
  NOR2_X1 u5_mult_82_U2870 ( .A1(u5_mult_82_n436), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__5_) );
  NOR2_X1 u5_mult_82_U2869 ( .A1(u5_mult_82_n434), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__6_) );
  NOR2_X1 u5_mult_82_U2868 ( .A1(u5_mult_82_n432), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__7_) );
  NOR2_X1 u5_mult_82_U2867 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__8_) );
  NOR2_X1 u5_mult_82_U2866 ( .A1(u5_mult_82_n428), .A2(u5_mult_82_n299), .ZN(
        u5_mult_82_ab_16__9_) );
  NOR2_X1 u5_mult_82_U2865 ( .A1(u5_mult_82_n480), .A2(u5_mult_82_n297), .ZN(
        u5_mult_82_ab_17__0_) );
  NOR2_X1 u5_mult_82_U2864 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n297), .ZN(
        u5_mult_82_ab_17__10_) );
  NOR2_X1 u5_mult_82_U2863 ( .A1(u5_mult_82_n426), .A2(u5_mult_82_n297), .ZN(
        u5_mult_82_ab_17__11_) );
  NOR2_X1 u5_mult_82_U2862 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n297), .ZN(
        u5_mult_82_ab_17__12_) );
  NOR2_X1 u5_mult_82_U2861 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n297), .ZN(
        u5_mult_82_ab_17__13_) );
  NOR2_X1 u5_mult_82_U2860 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n297), .ZN(
        u5_mult_82_ab_17__14_) );
  NOR2_X1 u5_mult_82_U2859 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n297), .ZN(
        u5_mult_82_ab_17__15_) );
  NOR2_X1 u5_mult_82_U2858 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n297), .ZN(
        u5_mult_82_ab_17__16_) );
  NOR2_X1 u5_mult_82_U2857 ( .A1(u5_mult_82_n409), .A2(u5_mult_82_n297), .ZN(
        u5_mult_82_ab_17__17_) );
  NOR2_X1 u5_mult_82_U2856 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n297), .ZN(
        u5_mult_82_ab_17__18_) );
  NOR2_X1 u5_mult_82_U2855 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n297), .ZN(
        u5_mult_82_ab_17__19_) );
  NOR2_X1 u5_mult_82_U2854 ( .A1(u5_mult_82_n443), .A2(u5_mult_82_n297), .ZN(
        u5_mult_82_ab_17__1_) );
  NOR2_X1 u5_mult_82_U2853 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n298), .ZN(
        u5_mult_82_ab_17__20_) );
  NOR2_X1 u5_mult_82_U2852 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n298), .ZN(
        u5_mult_82_ab_17__21_) );
  NOR2_X1 u5_mult_82_U2851 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n298), .ZN(
        u5_mult_82_ab_17__22_) );
  NOR2_X1 u5_mult_82_U2850 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n298), .ZN(
        u5_mult_82_ab_17__23_) );
  NOR2_X1 u5_mult_82_U2849 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n298), .ZN(
        u5_mult_82_ab_17__24_) );
  NOR2_X1 u5_mult_82_U2848 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n297), .ZN(
        u5_mult_82_ab_17__25_) );
  NOR2_X1 u5_mult_82_U2847 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n298), .ZN(
        u5_mult_82_ab_17__26_) );
  NOR2_X1 u5_mult_82_U2846 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n297), .ZN(
        u5_mult_82_ab_17__27_) );
  NOR2_X1 u5_mult_82_U2845 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n297), .ZN(
        u5_mult_82_ab_17__28_) );
  NOR2_X1 u5_mult_82_U2844 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n298), .ZN(
        u5_mult_82_ab_17__29_) );
  NOR2_X1 u5_mult_82_U2843 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n297), .ZN(
        u5_mult_82_ab_17__2_) );
  NOR2_X1 u5_mult_82_U2842 ( .A1(u5_mult_82_n384), .A2(u5_mult_82_n298), .ZN(
        u5_mult_82_ab_17__30_) );
  NOR2_X1 u5_mult_82_U2841 ( .A1(u5_mult_82_n382), .A2(u5_mult_82_n298), .ZN(
        u5_mult_82_ab_17__31_) );
  NOR2_X1 u5_mult_82_U2840 ( .A1(u5_mult_82_n380), .A2(u5_mult_82_n466), .ZN(
        u5_mult_82_ab_17__32_) );
  NOR2_X1 u5_mult_82_U2839 ( .A1(u5_mult_82_n378), .A2(u5_mult_82_n466), .ZN(
        u5_mult_82_ab_17__33_) );
  NOR2_X1 u5_mult_82_U2838 ( .A1(u5_mult_82_n376), .A2(u5_mult_82_n466), .ZN(
        u5_mult_82_ab_17__34_) );
  NOR2_X1 u5_mult_82_U2837 ( .A1(u5_mult_82_n374), .A2(u5_mult_82_n466), .ZN(
        u5_mult_82_ab_17__35_) );
  NOR2_X1 u5_mult_82_U2836 ( .A1(u5_mult_82_n474), .A2(u5_mult_82_n466), .ZN(
        u5_mult_82_ab_17__36_) );
  NOR2_X1 u5_mult_82_U2835 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n466), .ZN(
        u5_mult_82_ab_17__37_) );
  NOR2_X1 u5_mult_82_U2834 ( .A1(u5_mult_82_n367), .A2(u5_mult_82_n466), .ZN(
        u5_mult_82_ab_17__38_) );
  NOR2_X1 u5_mult_82_U2833 ( .A1(u5_mult_82_n366), .A2(u5_mult_82_n466), .ZN(
        u5_mult_82_ab_17__39_) );
  NOR2_X1 u5_mult_82_U2832 ( .A1(u5_mult_82_n441), .A2(u5_mult_82_n298), .ZN(
        u5_mult_82_ab_17__3_) );
  NOR2_X1 u5_mult_82_U2831 ( .A1(u5_mult_82_n364), .A2(u5_mult_82_n298), .ZN(
        u5_mult_82_ab_17__40_) );
  NOR2_X1 u5_mult_82_U2830 ( .A1(u5_mult_82_n362), .A2(u5_mult_82_n298), .ZN(
        u5_mult_82_ab_17__41_) );
  NOR2_X1 u5_mult_82_U2829 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n298), .ZN(
        u5_mult_82_ab_17__42_) );
  NOR2_X1 u5_mult_82_U2828 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n298), .ZN(
        u5_mult_82_ab_17__43_) );
  NOR2_X1 u5_mult_82_U2827 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n298), .ZN(
        u5_mult_82_ab_17__44_) );
  NOR2_X1 u5_mult_82_U2826 ( .A1(u5_mult_82_n352), .A2(u5_mult_82_n298), .ZN(
        u5_mult_82_ab_17__45_) );
  NOR2_X1 u5_mult_82_U2825 ( .A1(u5_mult_82_n350), .A2(u5_mult_82_n298), .ZN(
        u5_mult_82_ab_17__46_) );
  NOR2_X1 u5_mult_82_U2824 ( .A1(u5_mult_82_n348), .A2(u5_mult_82_n298), .ZN(
        u5_mult_82_ab_17__47_) );
  NOR2_X1 u5_mult_82_U2823 ( .A1(u5_mult_82_n346), .A2(u5_mult_82_n298), .ZN(
        u5_mult_82_ab_17__48_) );
  NOR2_X1 u5_mult_82_U2822 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n298), .ZN(
        u5_mult_82_ab_17__49_) );
  NOR2_X1 u5_mult_82_U2821 ( .A1(u5_mult_82_n438), .A2(u5_mult_82_n297), .ZN(
        u5_mult_82_ab_17__4_) );
  NOR2_X1 u5_mult_82_U2820 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n297), .ZN(
        u5_mult_82_ab_17__50_) );
  NOR2_X1 u5_mult_82_U2819 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n297), .ZN(
        u5_mult_82_ab_17__51_) );
  NOR2_X1 u5_mult_82_U2818 ( .A1(u5_mult_82_n336), .A2(u5_mult_82_n297), .ZN(
        u5_mult_82_ab_17__52_) );
  NOR2_X1 u5_mult_82_U2817 ( .A1(u5_mult_82_n436), .A2(u5_mult_82_n297), .ZN(
        u5_mult_82_ab_17__5_) );
  NOR2_X1 u5_mult_82_U2816 ( .A1(u5_mult_82_n434), .A2(u5_mult_82_n297), .ZN(
        u5_mult_82_ab_17__6_) );
  NOR2_X1 u5_mult_82_U2815 ( .A1(u5_mult_82_n432), .A2(u5_mult_82_n297), .ZN(
        u5_mult_82_ab_17__7_) );
  NOR2_X1 u5_mult_82_U2814 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n297), .ZN(
        u5_mult_82_ab_17__8_) );
  NOR2_X1 u5_mult_82_U2813 ( .A1(u5_mult_82_n428), .A2(u5_mult_82_n297), .ZN(
        u5_mult_82_ab_17__9_) );
  NOR2_X1 u5_mult_82_U2812 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n295), .ZN(
        u5_mult_82_ab_18__0_) );
  NOR2_X1 u5_mult_82_U2811 ( .A1(u5_mult_82_n477), .A2(u5_mult_82_n295), .ZN(
        u5_mult_82_ab_18__10_) );
  NOR2_X1 u5_mult_82_U2810 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n295), .ZN(
        u5_mult_82_ab_18__11_) );
  NOR2_X1 u5_mult_82_U2809 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n295), .ZN(
        u5_mult_82_ab_18__12_) );
  NOR2_X1 u5_mult_82_U2808 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n295), .ZN(
        u5_mult_82_ab_18__13_) );
  NOR2_X1 u5_mult_82_U2807 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n295), .ZN(
        u5_mult_82_ab_18__14_) );
  NOR2_X1 u5_mult_82_U2806 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n295), .ZN(
        u5_mult_82_ab_18__15_) );
  NOR2_X1 u5_mult_82_U2805 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n295), .ZN(
        u5_mult_82_ab_18__16_) );
  NOR2_X1 u5_mult_82_U2804 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n295), .ZN(
        u5_mult_82_ab_18__17_) );
  NOR2_X1 u5_mult_82_U2803 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n295), .ZN(
        u5_mult_82_ab_18__18_) );
  NOR2_X1 u5_mult_82_U2802 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n295), .ZN(
        u5_mult_82_ab_18__19_) );
  NOR2_X1 u5_mult_82_U2801 ( .A1(u5_mult_82_n443), .A2(u5_mult_82_n296), .ZN(
        u5_mult_82_ab_18__1_) );
  NOR2_X1 u5_mult_82_U2800 ( .A1(u5_mult_82_n475), .A2(u5_mult_82_n296), .ZN(
        u5_mult_82_ab_18__20_) );
  NOR2_X1 u5_mult_82_U2799 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n295), .ZN(
        u5_mult_82_ab_18__21_) );
  NOR2_X1 u5_mult_82_U2798 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n296), .ZN(
        u5_mult_82_ab_18__22_) );
  NOR2_X1 u5_mult_82_U2797 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n296), .ZN(
        u5_mult_82_ab_18__23_) );
  NOR2_X1 u5_mult_82_U2796 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n295), .ZN(
        u5_mult_82_ab_18__24_) );
  NOR2_X1 u5_mult_82_U2795 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n295), .ZN(
        u5_mult_82_ab_18__25_) );
  NOR2_X1 u5_mult_82_U2794 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n295), .ZN(
        u5_mult_82_ab_18__26_) );
  NOR2_X1 u5_mult_82_U2793 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n295), .ZN(
        u5_mult_82_ab_18__27_) );
  NOR2_X1 u5_mult_82_U2792 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n296), .ZN(
        u5_mult_82_ab_18__28_) );
  NOR2_X1 u5_mult_82_U2791 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n296), .ZN(
        u5_mult_82_ab_18__29_) );
  NOR2_X1 u5_mult_82_U2790 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n295), .ZN(
        u5_mult_82_ab_18__2_) );
  NOR2_X1 u5_mult_82_U2789 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n296), .ZN(
        u5_mult_82_ab_18__30_) );
  NOR2_X1 u5_mult_82_U2788 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n296), .ZN(
        u5_mult_82_ab_18__31_) );
  NOR2_X1 u5_mult_82_U2787 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n465), .ZN(
        u5_mult_82_ab_18__32_) );
  NOR2_X1 u5_mult_82_U2786 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n465), .ZN(
        u5_mult_82_ab_18__33_) );
  NOR2_X1 u5_mult_82_U2785 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n465), .ZN(
        u5_mult_82_ab_18__34_) );
  NOR2_X1 u5_mult_82_U2784 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n465), .ZN(
        u5_mult_82_ab_18__35_) );
  NOR2_X1 u5_mult_82_U2783 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n465), .ZN(
        u5_mult_82_ab_18__36_) );
  NOR2_X1 u5_mult_82_U2782 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n465), .ZN(
        u5_mult_82_ab_18__37_) );
  NOR2_X1 u5_mult_82_U2781 ( .A1(u5_mult_82_n367), .A2(u5_mult_82_n465), .ZN(
        u5_mult_82_ab_18__38_) );
  NOR2_X1 u5_mult_82_U2780 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n295), .ZN(
        u5_mult_82_ab_18__39_) );
  NOR2_X1 u5_mult_82_U2779 ( .A1(u5_mult_82_n441), .A2(u5_mult_82_n296), .ZN(
        u5_mult_82_ab_18__3_) );
  NOR2_X1 u5_mult_82_U2778 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n296), .ZN(
        u5_mult_82_ab_18__40_) );
  NOR2_X1 u5_mult_82_U2777 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n296), .ZN(
        u5_mult_82_ab_18__41_) );
  NOR2_X1 u5_mult_82_U2776 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n296), .ZN(
        u5_mult_82_ab_18__42_) );
  NOR2_X1 u5_mult_82_U2775 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n296), .ZN(
        u5_mult_82_ab_18__43_) );
  NOR2_X1 u5_mult_82_U2774 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n296), .ZN(
        u5_mult_82_ab_18__44_) );
  NOR2_X1 u5_mult_82_U2773 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n296), .ZN(
        u5_mult_82_ab_18__45_) );
  NOR2_X1 u5_mult_82_U2772 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n296), .ZN(
        u5_mult_82_ab_18__46_) );
  NOR2_X1 u5_mult_82_U2771 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n296), .ZN(
        u5_mult_82_ab_18__47_) );
  NOR2_X1 u5_mult_82_U2770 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n296), .ZN(
        u5_mult_82_ab_18__48_) );
  NOR2_X1 u5_mult_82_U2769 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n296), .ZN(
        u5_mult_82_ab_18__49_) );
  NOR2_X1 u5_mult_82_U2768 ( .A1(u5_mult_82_n438), .A2(u5_mult_82_n295), .ZN(
        u5_mult_82_ab_18__4_) );
  NOR2_X1 u5_mult_82_U2767 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n295), .ZN(
        u5_mult_82_ab_18__50_) );
  NOR2_X1 u5_mult_82_U2766 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n295), .ZN(
        u5_mult_82_ab_18__51_) );
  NOR2_X1 u5_mult_82_U2765 ( .A1(u5_mult_82_n336), .A2(u5_mult_82_n295), .ZN(
        u5_mult_82_ab_18__52_) );
  NOR2_X1 u5_mult_82_U2764 ( .A1(u5_mult_82_n436), .A2(u5_mult_82_n295), .ZN(
        u5_mult_82_ab_18__5_) );
  NOR2_X1 u5_mult_82_U2763 ( .A1(u5_mult_82_n434), .A2(u5_mult_82_n295), .ZN(
        u5_mult_82_ab_18__6_) );
  NOR2_X1 u5_mult_82_U2762 ( .A1(u5_mult_82_n432), .A2(u5_mult_82_n295), .ZN(
        u5_mult_82_ab_18__7_) );
  NOR2_X1 u5_mult_82_U2761 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n295), .ZN(
        u5_mult_82_ab_18__8_) );
  NOR2_X1 u5_mult_82_U2760 ( .A1(u5_mult_82_n428), .A2(u5_mult_82_n295), .ZN(
        u5_mult_82_ab_18__9_) );
  NOR2_X1 u5_mult_82_U2759 ( .A1(u5_mult_82_n480), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__0_) );
  NOR2_X1 u5_mult_82_U2758 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__10_) );
  NOR2_X1 u5_mult_82_U2757 ( .A1(u5_mult_82_n426), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__11_) );
  NOR2_X1 u5_mult_82_U2756 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__12_) );
  NOR2_X1 u5_mult_82_U2755 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__13_) );
  NOR2_X1 u5_mult_82_U2754 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__14_) );
  NOR2_X1 u5_mult_82_U2753 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__15_) );
  NOR2_X1 u5_mult_82_U2752 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__16_) );
  NOR2_X1 u5_mult_82_U2751 ( .A1(u5_mult_82_n409), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__17_) );
  NOR2_X1 u5_mult_82_U2750 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__18_) );
  NOR2_X1 u5_mult_82_U2749 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__19_) );
  NOR2_X1 u5_mult_82_U2748 ( .A1(u5_mult_82_n443), .A2(u5_mult_82_n293), .ZN(
        u5_mult_82_ab_19__1_) );
  NOR2_X1 u5_mult_82_U2747 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n293), .ZN(
        u5_mult_82_ab_19__20_) );
  NOR2_X1 u5_mult_82_U2746 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n293), .ZN(
        u5_mult_82_ab_19__21_) );
  NOR2_X1 u5_mult_82_U2745 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n293), .ZN(
        u5_mult_82_ab_19__22_) );
  NOR2_X1 u5_mult_82_U2744 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n293), .ZN(
        u5_mult_82_ab_19__23_) );
  NOR2_X1 u5_mult_82_U2743 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n293), .ZN(
        u5_mult_82_ab_19__24_) );
  NOR2_X1 u5_mult_82_U2742 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__25_) );
  NOR2_X1 u5_mult_82_U2741 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__26_) );
  NOR2_X1 u5_mult_82_U2740 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__27_) );
  NOR2_X1 u5_mult_82_U2739 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__28_) );
  NOR2_X1 u5_mult_82_U2738 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__29_) );
  NOR2_X1 u5_mult_82_U2737 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n293), .ZN(
        u5_mult_82_ab_19__2_) );
  NOR2_X1 u5_mult_82_U2736 ( .A1(u5_mult_82_n384), .A2(u5_mult_82_n293), .ZN(
        u5_mult_82_ab_19__30_) );
  NOR2_X1 u5_mult_82_U2735 ( .A1(u5_mult_82_n382), .A2(u5_mult_82_n293), .ZN(
        u5_mult_82_ab_19__31_) );
  NOR2_X1 u5_mult_82_U2734 ( .A1(u5_mult_82_n380), .A2(u5_mult_82_n293), .ZN(
        u5_mult_82_ab_19__32_) );
  NOR2_X1 u5_mult_82_U2733 ( .A1(u5_mult_82_n378), .A2(u5_mult_82_n293), .ZN(
        u5_mult_82_ab_19__33_) );
  NOR2_X1 u5_mult_82_U2732 ( .A1(u5_mult_82_n376), .A2(u5_mult_82_n293), .ZN(
        u5_mult_82_ab_19__34_) );
  NOR2_X1 u5_mult_82_U2731 ( .A1(u5_mult_82_n374), .A2(u5_mult_82_n293), .ZN(
        u5_mult_82_ab_19__35_) );
  NOR2_X1 u5_mult_82_U2730 ( .A1(u5_mult_82_n474), .A2(u5_mult_82_n293), .ZN(
        u5_mult_82_ab_19__36_) );
  NOR2_X1 u5_mult_82_U2729 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n293), .ZN(
        u5_mult_82_ab_19__37_) );
  NOR2_X1 u5_mult_82_U2728 ( .A1(u5_mult_82_n367), .A2(u5_mult_82_n293), .ZN(
        u5_mult_82_ab_19__38_) );
  NOR2_X1 u5_mult_82_U2727 ( .A1(u5_mult_82_n366), .A2(u5_mult_82_n293), .ZN(
        u5_mult_82_ab_19__39_) );
  NOR2_X1 u5_mult_82_U2726 ( .A1(u5_mult_82_n441), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__3_) );
  NOR2_X1 u5_mult_82_U2725 ( .A1(u5_mult_82_n364), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__40_) );
  NOR2_X1 u5_mult_82_U2724 ( .A1(u5_mult_82_n362), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__41_) );
  NOR2_X1 u5_mult_82_U2723 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__42_) );
  NOR2_X1 u5_mult_82_U2722 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__43_) );
  NOR2_X1 u5_mult_82_U2721 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__44_) );
  NOR2_X1 u5_mult_82_U2720 ( .A1(u5_mult_82_n352), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__45_) );
  NOR2_X1 u5_mult_82_U2719 ( .A1(u5_mult_82_n350), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__46_) );
  NOR2_X1 u5_mult_82_U2718 ( .A1(u5_mult_82_n348), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__47_) );
  NOR2_X1 u5_mult_82_U2717 ( .A1(u5_mult_82_n346), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__48_) );
  NOR2_X1 u5_mult_82_U2716 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__49_) );
  NOR2_X1 u5_mult_82_U2715 ( .A1(u5_mult_82_n438), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__4_) );
  NOR2_X1 u5_mult_82_U2714 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__50_) );
  NOR2_X1 u5_mult_82_U2713 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__51_) );
  NOR2_X1 u5_mult_82_U2712 ( .A1(u5_mult_82_n336), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__52_) );
  NOR2_X1 u5_mult_82_U2711 ( .A1(u5_mult_82_n436), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__5_) );
  NOR2_X1 u5_mult_82_U2710 ( .A1(u5_mult_82_n434), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__6_) );
  NOR2_X1 u5_mult_82_U2709 ( .A1(u5_mult_82_n432), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__7_) );
  NOR2_X1 u5_mult_82_U2708 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__8_) );
  NOR2_X1 u5_mult_82_U2707 ( .A1(u5_mult_82_n428), .A2(u5_mult_82_n294), .ZN(
        u5_mult_82_ab_19__9_) );
  NOR2_X1 u5_mult_82_U2706 ( .A1(u5_mult_82_n480), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__0_) );
  NOR2_X1 u5_mult_82_U2705 ( .A1(u5_mult_82_n477), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__10_) );
  NOR2_X1 u5_mult_82_U2704 ( .A1(u5_mult_82_n426), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__11_) );
  NOR2_X1 u5_mult_82_U2703 ( .A1(u5_mult_82_n422), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__12_) );
  NOR2_X1 u5_mult_82_U2702 ( .A1(u5_mult_82_n419), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__13_) );
  NOR2_X1 u5_mult_82_U2701 ( .A1(u5_mult_82_n416), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__14_) );
  NOR2_X1 u5_mult_82_U2700 ( .A1(u5_mult_82_n413), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__15_) );
  NOR2_X1 u5_mult_82_U2699 ( .A1(u5_mult_82_n410), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__16_) );
  NOR2_X1 u5_mult_82_U2698 ( .A1(u5_mult_82_n409), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__17_) );
  NOR2_X1 u5_mult_82_U2697 ( .A1(u5_mult_82_n476), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__18_) );
  NOR2_X1 u5_mult_82_U2696 ( .A1(u5_mult_82_n404), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__19_) );
  NOR2_X1 u5_mult_82_U2695 ( .A1(u5_mult_82_n445), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__1_) );
  NOR2_X1 u5_mult_82_U2694 ( .A1(u5_mult_82_n475), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__20_) );
  NOR2_X1 u5_mult_82_U2693 ( .A1(u5_mult_82_n402), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__21_) );
  NOR2_X1 u5_mult_82_U2692 ( .A1(u5_mult_82_n400), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__22_) );
  NOR2_X1 u5_mult_82_U2691 ( .A1(u5_mult_82_n398), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__23_) );
  NOR2_X1 u5_mult_82_U2690 ( .A1(u5_mult_82_n396), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__24_) );
  NOR2_X1 u5_mult_82_U2689 ( .A1(u5_mult_82_n394), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__25_) );
  NOR2_X1 u5_mult_82_U2688 ( .A1(u5_mult_82_n392), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__26_) );
  NOR2_X1 u5_mult_82_U2687 ( .A1(u5_mult_82_n390), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__27_) );
  NOR2_X1 u5_mult_82_U2686 ( .A1(u5_mult_82_n387), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__28_) );
  NOR2_X1 u5_mult_82_U2685 ( .A1(u5_mult_82_n386), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__29_) );
  NOR2_X1 u5_mult_82_U2684 ( .A1(u5_mult_82_n442), .A2(u5_mult_82_n331), .ZN(
        u5_mult_82_ab_1__2_) );
  NOR2_X1 u5_mult_82_U2683 ( .A1(u5_mult_82_n384), .A2(u5_mult_82_n331), .ZN(
        u5_mult_82_ab_1__30_) );
  NOR2_X1 u5_mult_82_U2682 ( .A1(u5_mult_82_n382), .A2(u5_mult_82_n331), .ZN(
        u5_mult_82_ab_1__31_) );
  NOR2_X1 u5_mult_82_U2681 ( .A1(u5_mult_82_n380), .A2(u5_mult_82_n331), .ZN(
        u5_mult_82_ab_1__32_) );
  NOR2_X1 u5_mult_82_U2680 ( .A1(u5_mult_82_n378), .A2(u5_mult_82_n331), .ZN(
        u5_mult_82_ab_1__33_) );
  NOR2_X1 u5_mult_82_U2679 ( .A1(u5_mult_82_n376), .A2(u5_mult_82_n331), .ZN(
        u5_mult_82_ab_1__34_) );
  NOR2_X1 u5_mult_82_U2678 ( .A1(u5_mult_82_n374), .A2(u5_mult_82_n331), .ZN(
        u5_mult_82_ab_1__35_) );
  NOR2_X1 u5_mult_82_U2677 ( .A1(u5_mult_82_n474), .A2(u5_mult_82_n331), .ZN(
        u5_mult_82_ab_1__36_) );
  NOR2_X1 u5_mult_82_U2676 ( .A1(u5_mult_82_n370), .A2(u5_mult_82_n331), .ZN(
        u5_mult_82_ab_1__37_) );
  NOR2_X1 u5_mult_82_U2675 ( .A1(u5_mult_82_n368), .A2(u5_mult_82_n331), .ZN(
        u5_mult_82_ab_1__38_) );
  NOR2_X1 u5_mult_82_U2674 ( .A1(u5_mult_82_n366), .A2(u5_mult_82_n331), .ZN(
        u5_mult_82_ab_1__39_) );
  NOR2_X1 u5_mult_82_U2673 ( .A1(u5_mult_82_n440), .A2(u5_mult_82_n332), .ZN(
        u5_mult_82_ab_1__3_) );
  NOR2_X1 u5_mult_82_U2672 ( .A1(u5_mult_82_n364), .A2(u5_mult_82_n332), .ZN(
        u5_mult_82_ab_1__40_) );
  NOR2_X1 u5_mult_82_U2671 ( .A1(u5_mult_82_n362), .A2(u5_mult_82_n332), .ZN(
        u5_mult_82_ab_1__41_) );
  NOR2_X1 u5_mult_82_U2670 ( .A1(u5_mult_82_n358), .A2(u5_mult_82_n332), .ZN(
        u5_mult_82_ab_1__42_) );
  NOR2_X1 u5_mult_82_U2669 ( .A1(u5_mult_82_n356), .A2(u5_mult_82_n332), .ZN(
        u5_mult_82_ab_1__43_) );
  NOR2_X1 u5_mult_82_U2668 ( .A1(u5_mult_82_n353), .A2(u5_mult_82_n332), .ZN(
        u5_mult_82_ab_1__44_) );
  NOR2_X1 u5_mult_82_U2667 ( .A1(u5_mult_82_n352), .A2(u5_mult_82_n332), .ZN(
        u5_mult_82_ab_1__45_) );
  NOR2_X1 u5_mult_82_U2666 ( .A1(u5_mult_82_n350), .A2(u5_mult_82_n332), .ZN(
        u5_mult_82_ab_1__46_) );
  NOR2_X1 u5_mult_82_U2665 ( .A1(u5_mult_82_n348), .A2(u5_mult_82_n332), .ZN(
        u5_mult_82_ab_1__47_) );
  NOR2_X1 u5_mult_82_U2664 ( .A1(u5_mult_82_n346), .A2(u5_mult_82_n332), .ZN(
        u5_mult_82_ab_1__48_) );
  NOR2_X1 u5_mult_82_U2663 ( .A1(u5_mult_82_n343), .A2(u5_mult_82_n332), .ZN(
        u5_mult_82_ab_1__49_) );
  NOR2_X1 u5_mult_82_U2662 ( .A1(u5_mult_82_n438), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__4_) );
  NOR2_X1 u5_mult_82_U2661 ( .A1(u5_mult_82_n342), .A2(u5_mult_82_n332), .ZN(
        u5_mult_82_ab_1__50_) );
  NOR2_X1 u5_mult_82_U2660 ( .A1(u5_mult_82_n340), .A2(u5_mult_82_n331), .ZN(
        u5_mult_82_ab_1__51_) );
  NOR2_X1 u5_mult_82_U2659 ( .A1(u5_mult_82_n336), .A2(u5_mult_82_n331), .ZN(
        u5_mult_82_ab_1__52_) );
  NOR2_X1 u5_mult_82_U2658 ( .A1(u5_mult_82_n436), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__5_) );
  NOR2_X1 u5_mult_82_U2657 ( .A1(u5_mult_82_n434), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__6_) );
  NOR2_X1 u5_mult_82_U2656 ( .A1(u5_mult_82_n432), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__7_) );
  NOR2_X1 u5_mult_82_U2655 ( .A1(u5_mult_82_n430), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__8_) );
  NOR2_X1 u5_mult_82_U2654 ( .A1(u5_mult_82_n428), .A2(u5_mult_82_n330), .ZN(
        u5_mult_82_ab_1__9_) );
  NOR2_X1 u5_mult_82_U2653 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__0_) );
  NOR2_X1 u5_mult_82_U2652 ( .A1(u5_mult_82_n477), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__10_) );
  NOR2_X1 u5_mult_82_U2651 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__11_) );
  NOR2_X1 u5_mult_82_U2650 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__12_) );
  NOR2_X1 u5_mult_82_U2649 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__13_) );
  NOR2_X1 u5_mult_82_U2648 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__14_) );
  NOR2_X1 u5_mult_82_U2647 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__15_) );
  NOR2_X1 u5_mult_82_U2646 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__16_) );
  NOR2_X1 u5_mult_82_U2645 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__17_) );
  NOR2_X1 u5_mult_82_U2644 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__18_) );
  NOR2_X1 u5_mult_82_U2643 ( .A1(u5_mult_82_n404), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__19_) );
  NOR2_X1 u5_mult_82_U2642 ( .A1(u5_mult_82_n443), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__1_) );
  NOR2_X1 u5_mult_82_U2641 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__20_) );
  NOR2_X1 u5_mult_82_U2640 ( .A1(u5_mult_82_n402), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__21_) );
  NOR2_X1 u5_mult_82_U2639 ( .A1(u5_mult_82_n400), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__22_) );
  NOR2_X1 u5_mult_82_U2638 ( .A1(u5_mult_82_n398), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__23_) );
  NOR2_X1 u5_mult_82_U2637 ( .A1(u5_mult_82_n396), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__24_) );
  NOR2_X1 u5_mult_82_U2636 ( .A1(u5_mult_82_n394), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__25_) );
  NOR2_X1 u5_mult_82_U2635 ( .A1(u5_mult_82_n392), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__26_) );
  NOR2_X1 u5_mult_82_U2634 ( .A1(u5_mult_82_n390), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__27_) );
  NOR2_X1 u5_mult_82_U2633 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__28_) );
  NOR2_X1 u5_mult_82_U2632 ( .A1(u5_mult_82_n386), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__29_) );
  NOR2_X1 u5_mult_82_U2631 ( .A1(u5_mult_82_n442), .A2(u5_mult_82_n464), .ZN(
        u5_mult_82_ab_20__2_) );
  NOR2_X1 u5_mult_82_U2630 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n464), .ZN(
        u5_mult_82_ab_20__30_) );
  NOR2_X1 u5_mult_82_U2629 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n464), .ZN(
        u5_mult_82_ab_20__31_) );
  NOR2_X1 u5_mult_82_U2628 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n464), .ZN(
        u5_mult_82_ab_20__32_) );
  NOR2_X1 u5_mult_82_U2627 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n464), .ZN(
        u5_mult_82_ab_20__33_) );
  NOR2_X1 u5_mult_82_U2626 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n464), .ZN(
        u5_mult_82_ab_20__34_) );
  NOR2_X1 u5_mult_82_U2625 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n464), .ZN(
        u5_mult_82_ab_20__35_) );
  NOR2_X1 u5_mult_82_U2624 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n464), .ZN(
        u5_mult_82_ab_20__36_) );
  NOR2_X1 u5_mult_82_U2623 ( .A1(u5_mult_82_n370), .A2(u5_mult_82_n464), .ZN(
        u5_mult_82_ab_20__37_) );
  NOR2_X1 u5_mult_82_U2622 ( .A1(u5_mult_82_n368), .A2(u5_mult_82_n464), .ZN(
        u5_mult_82_ab_20__38_) );
  NOR2_X1 u5_mult_82_U2621 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n464), .ZN(
        u5_mult_82_ab_20__39_) );
  NOR2_X1 u5_mult_82_U2620 ( .A1(u5_mult_82_n440), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__3_) );
  NOR2_X1 u5_mult_82_U2619 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__40_) );
  NOR2_X1 u5_mult_82_U2618 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__41_) );
  NOR2_X1 u5_mult_82_U2617 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__42_) );
  NOR2_X1 u5_mult_82_U2616 ( .A1(u5_mult_82_n356), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__43_) );
  NOR2_X1 u5_mult_82_U2615 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__44_) );
  NOR2_X1 u5_mult_82_U2614 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__45_) );
  NOR2_X1 u5_mult_82_U2613 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__46_) );
  NOR2_X1 u5_mult_82_U2612 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__47_) );
  NOR2_X1 u5_mult_82_U2611 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__48_) );
  NOR2_X1 u5_mult_82_U2610 ( .A1(u5_mult_82_n343), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__49_) );
  NOR2_X1 u5_mult_82_U2609 ( .A1(u5_mult_82_n438), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__4_) );
  NOR2_X1 u5_mult_82_U2608 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__50_) );
  NOR2_X1 u5_mult_82_U2607 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__51_) );
  NOR2_X1 u5_mult_82_U2606 ( .A1(u5_mult_82_n336), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__52_) );
  NOR2_X1 u5_mult_82_U2605 ( .A1(u5_mult_82_n436), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__5_) );
  NOR2_X1 u5_mult_82_U2604 ( .A1(u5_mult_82_n434), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__6_) );
  NOR2_X1 u5_mult_82_U2603 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__7_) );
  NOR2_X1 u5_mult_82_U2602 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__8_) );
  NOR2_X1 u5_mult_82_U2601 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n292), .ZN(
        u5_mult_82_ab_20__9_) );
  NOR2_X1 u5_mult_82_U2600 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__0_) );
  NOR2_X1 u5_mult_82_U2599 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__10_) );
  NOR2_X1 u5_mult_82_U2598 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__11_) );
  NOR2_X1 u5_mult_82_U2597 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__12_) );
  NOR2_X1 u5_mult_82_U2596 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__13_) );
  NOR2_X1 u5_mult_82_U2595 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__14_) );
  NOR2_X1 u5_mult_82_U2594 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__15_) );
  NOR2_X1 u5_mult_82_U2593 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__16_) );
  NOR2_X1 u5_mult_82_U2592 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__17_) );
  NOR2_X1 u5_mult_82_U2591 ( .A1(u5_mult_82_n406), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__18_) );
  NOR2_X1 u5_mult_82_U2590 ( .A1(u5_mult_82_n404), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__19_) );
  NOR2_X1 u5_mult_82_U2589 ( .A1(u5_mult_82_n443), .A2(u5_mult_82_n463), .ZN(
        u5_mult_82_ab_21__1_) );
  NOR2_X1 u5_mult_82_U2588 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n463), .ZN(
        u5_mult_82_ab_21__20_) );
  NOR2_X1 u5_mult_82_U2587 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n463), .ZN(
        u5_mult_82_ab_21__21_) );
  NOR2_X1 u5_mult_82_U2586 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__22_) );
  NOR2_X1 u5_mult_82_U2585 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n290), .ZN(
        u5_mult_82_ab_21__23_) );
  NOR2_X1 u5_mult_82_U2584 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n290), .ZN(
        u5_mult_82_ab_21__24_) );
  NOR2_X1 u5_mult_82_U2583 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n290), .ZN(
        u5_mult_82_ab_21__25_) );
  NOR2_X1 u5_mult_82_U2582 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n290), .ZN(
        u5_mult_82_ab_21__26_) );
  NOR2_X1 u5_mult_82_U2581 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__27_) );
  NOR2_X1 u5_mult_82_U2580 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n290), .ZN(
        u5_mult_82_ab_21__28_) );
  NOR2_X1 u5_mult_82_U2579 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n290), .ZN(
        u5_mult_82_ab_21__29_) );
  NOR2_X1 u5_mult_82_U2578 ( .A1(u5_mult_82_n442), .A2(u5_mult_82_n290), .ZN(
        u5_mult_82_ab_21__2_) );
  NOR2_X1 u5_mult_82_U2577 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n290), .ZN(
        u5_mult_82_ab_21__30_) );
  NOR2_X1 u5_mult_82_U2576 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n290), .ZN(
        u5_mult_82_ab_21__31_) );
  NOR2_X1 u5_mult_82_U2575 ( .A1(u5_mult_82_n380), .A2(u5_mult_82_n290), .ZN(
        u5_mult_82_ab_21__32_) );
  NOR2_X1 u5_mult_82_U2574 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n290), .ZN(
        u5_mult_82_ab_21__33_) );
  NOR2_X1 u5_mult_82_U2573 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n290), .ZN(
        u5_mult_82_ab_21__34_) );
  NOR2_X1 u5_mult_82_U2572 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n290), .ZN(
        u5_mult_82_ab_21__35_) );
  NOR2_X1 u5_mult_82_U2571 ( .A1(u5_mult_82_n474), .A2(u5_mult_82_n290), .ZN(
        u5_mult_82_ab_21__36_) );
  NOR2_X1 u5_mult_82_U2570 ( .A1(u5_mult_82_n370), .A2(u5_mult_82_n290), .ZN(
        u5_mult_82_ab_21__37_) );
  NOR2_X1 u5_mult_82_U2569 ( .A1(u5_mult_82_n368), .A2(u5_mult_82_n290), .ZN(
        u5_mult_82_ab_21__38_) );
  NOR2_X1 u5_mult_82_U2568 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n290), .ZN(
        u5_mult_82_ab_21__39_) );
  NOR2_X1 u5_mult_82_U2567 ( .A1(u5_mult_82_n440), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__3_) );
  NOR2_X1 u5_mult_82_U2566 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__40_) );
  NOR2_X1 u5_mult_82_U2565 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__41_) );
  NOR2_X1 u5_mult_82_U2564 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__42_) );
  NOR2_X1 u5_mult_82_U2563 ( .A1(u5_mult_82_n356), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__43_) );
  NOR2_X1 u5_mult_82_U2562 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__44_) );
  NOR2_X1 u5_mult_82_U2561 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__45_) );
  NOR2_X1 u5_mult_82_U2560 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__46_) );
  NOR2_X1 u5_mult_82_U2559 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__47_) );
  NOR2_X1 u5_mult_82_U2558 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__48_) );
  NOR2_X1 u5_mult_82_U2557 ( .A1(u5_mult_82_n343), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__49_) );
  NOR2_X1 u5_mult_82_U2556 ( .A1(u5_mult_82_n438), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__4_) );
  NOR2_X1 u5_mult_82_U2555 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__50_) );
  NOR2_X1 u5_mult_82_U2554 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__51_) );
  NOR2_X1 u5_mult_82_U2553 ( .A1(u5_mult_82_n336), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__52_) );
  NOR2_X1 u5_mult_82_U2552 ( .A1(u5_mult_82_n436), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__5_) );
  NOR2_X1 u5_mult_82_U2551 ( .A1(u5_mult_82_n434), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__6_) );
  NOR2_X1 u5_mult_82_U2550 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__7_) );
  NOR2_X1 u5_mult_82_U2549 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__8_) );
  NOR2_X1 u5_mult_82_U2548 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n291), .ZN(
        u5_mult_82_ab_21__9_) );
  NOR2_X1 u5_mult_82_U2547 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__0_) );
  NOR2_X1 u5_mult_82_U2546 ( .A1(u5_mult_82_n477), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__10_) );
  NOR2_X1 u5_mult_82_U2545 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__11_) );
  NOR2_X1 u5_mult_82_U2544 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__12_) );
  NOR2_X1 u5_mult_82_U2543 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__13_) );
  NOR2_X1 u5_mult_82_U2542 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__14_) );
  NOR2_X1 u5_mult_82_U2541 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__15_) );
  NOR2_X1 u5_mult_82_U2540 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__16_) );
  NOR2_X1 u5_mult_82_U2539 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__17_) );
  NOR2_X1 u5_mult_82_U2538 ( .A1(u5_mult_82_n406), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__18_) );
  NOR2_X1 u5_mult_82_U2537 ( .A1(u5_mult_82_n404), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__19_) );
  NOR2_X1 u5_mult_82_U2536 ( .A1(u5_mult_82_n443), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__1_) );
  NOR2_X1 u5_mult_82_U2535 ( .A1(u5_mult_82_n475), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__20_) );
  NOR2_X1 u5_mult_82_U2534 ( .A1(u5_mult_82_n402), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__21_) );
  NOR2_X1 u5_mult_82_U2533 ( .A1(u5_mult_82_n400), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__22_) );
  NOR2_X1 u5_mult_82_U2532 ( .A1(u5_mult_82_n398), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__23_) );
  NOR2_X1 u5_mult_82_U2531 ( .A1(u5_mult_82_n396), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__24_) );
  NOR2_X1 u5_mult_82_U2530 ( .A1(u5_mult_82_n394), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__25_) );
  NOR2_X1 u5_mult_82_U2529 ( .A1(u5_mult_82_n392), .A2(u5_mult_82_n288), .ZN(
        u5_mult_82_ab_22__26_) );
  NOR2_X1 u5_mult_82_U2528 ( .A1(u5_mult_82_n390), .A2(u5_mult_82_n288), .ZN(
        u5_mult_82_ab_22__27_) );
  NOR2_X1 u5_mult_82_U2527 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n288), .ZN(
        u5_mult_82_ab_22__28_) );
  NOR2_X1 u5_mult_82_U2526 ( .A1(u5_mult_82_n386), .A2(u5_mult_82_n288), .ZN(
        u5_mult_82_ab_22__29_) );
  NOR2_X1 u5_mult_82_U2525 ( .A1(u5_mult_82_n442), .A2(u5_mult_82_n288), .ZN(
        u5_mult_82_ab_22__2_) );
  NOR2_X1 u5_mult_82_U2524 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n288), .ZN(
        u5_mult_82_ab_22__30_) );
  NOR2_X1 u5_mult_82_U2523 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n288), .ZN(
        u5_mult_82_ab_22__31_) );
  NOR2_X1 u5_mult_82_U2522 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n288), .ZN(
        u5_mult_82_ab_22__32_) );
  NOR2_X1 u5_mult_82_U2521 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n288), .ZN(
        u5_mult_82_ab_22__33_) );
  NOR2_X1 u5_mult_82_U2520 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n288), .ZN(
        u5_mult_82_ab_22__34_) );
  NOR2_X1 u5_mult_82_U2519 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n288), .ZN(
        u5_mult_82_ab_22__35_) );
  NOR2_X1 u5_mult_82_U2518 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n288), .ZN(
        u5_mult_82_ab_22__36_) );
  NOR2_X1 u5_mult_82_U2517 ( .A1(u5_mult_82_n370), .A2(u5_mult_82_n288), .ZN(
        u5_mult_82_ab_22__37_) );
  NOR2_X1 u5_mult_82_U2516 ( .A1(u5_mult_82_n369), .A2(u5_mult_82_n288), .ZN(
        u5_mult_82_ab_22__38_) );
  NOR2_X1 u5_mult_82_U2515 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n288), .ZN(
        u5_mult_82_ab_22__39_) );
  NOR2_X1 u5_mult_82_U2514 ( .A1(u5_mult_82_n440), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__3_) );
  NOR2_X1 u5_mult_82_U2513 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__40_) );
  NOR2_X1 u5_mult_82_U2512 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__41_) );
  NOR2_X1 u5_mult_82_U2511 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__42_) );
  NOR2_X1 u5_mult_82_U2510 ( .A1(u5_mult_82_n356), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__43_) );
  NOR2_X1 u5_mult_82_U2509 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__44_) );
  NOR2_X1 u5_mult_82_U2508 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__45_) );
  NOR2_X1 u5_mult_82_U2507 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__46_) );
  NOR2_X1 u5_mult_82_U2506 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__47_) );
  NOR2_X1 u5_mult_82_U2505 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__48_) );
  NOR2_X1 u5_mult_82_U2504 ( .A1(u5_mult_82_n343), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__49_) );
  NOR2_X1 u5_mult_82_U2503 ( .A1(u5_mult_82_n438), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__4_) );
  NOR2_X1 u5_mult_82_U2502 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__50_) );
  NOR2_X1 u5_mult_82_U2501 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__51_) );
  NOR2_X1 u5_mult_82_U2500 ( .A1(u5_mult_82_n336), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__52_) );
  NOR2_X1 u5_mult_82_U2499 ( .A1(u5_mult_82_n436), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__5_) );
  NOR2_X1 u5_mult_82_U2498 ( .A1(u5_mult_82_n434), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__6_) );
  NOR2_X1 u5_mult_82_U2497 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__7_) );
  NOR2_X1 u5_mult_82_U2496 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__8_) );
  NOR2_X1 u5_mult_82_U2495 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n289), .ZN(
        u5_mult_82_ab_22__9_) );
  NOR2_X1 u5_mult_82_U2494 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__0_) );
  NOR2_X1 u5_mult_82_U2493 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__10_) );
  NOR2_X1 u5_mult_82_U2492 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__11_) );
  NOR2_X1 u5_mult_82_U2491 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__12_) );
  NOR2_X1 u5_mult_82_U2490 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__13_) );
  NOR2_X1 u5_mult_82_U2489 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__14_) );
  NOR2_X1 u5_mult_82_U2488 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__15_) );
  NOR2_X1 u5_mult_82_U2487 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__16_) );
  NOR2_X1 u5_mult_82_U2486 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__17_) );
  NOR2_X1 u5_mult_82_U2485 ( .A1(u5_mult_82_n406), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__18_) );
  NOR2_X1 u5_mult_82_U2484 ( .A1(u5_mult_82_n404), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__19_) );
  NOR2_X1 u5_mult_82_U2483 ( .A1(u5_mult_82_n443), .A2(u5_mult_82_n286), .ZN(
        u5_mult_82_ab_23__1_) );
  NOR2_X1 u5_mult_82_U2482 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__20_) );
  NOR2_X1 u5_mult_82_U2481 ( .A1(u5_mult_82_n402), .A2(u5_mult_82_n286), .ZN(
        u5_mult_82_ab_23__21_) );
  NOR2_X1 u5_mult_82_U2480 ( .A1(u5_mult_82_n400), .A2(u5_mult_82_n286), .ZN(
        u5_mult_82_ab_23__22_) );
  NOR2_X1 u5_mult_82_U2479 ( .A1(u5_mult_82_n398), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__23_) );
  NOR2_X1 u5_mult_82_U2478 ( .A1(u5_mult_82_n396), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__24_) );
  NOR2_X1 u5_mult_82_U2477 ( .A1(u5_mult_82_n394), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__25_) );
  NOR2_X1 u5_mult_82_U2476 ( .A1(u5_mult_82_n392), .A2(u5_mult_82_n286), .ZN(
        u5_mult_82_ab_23__26_) );
  NOR2_X1 u5_mult_82_U2475 ( .A1(u5_mult_82_n390), .A2(u5_mult_82_n286), .ZN(
        u5_mult_82_ab_23__27_) );
  NOR2_X1 u5_mult_82_U2474 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n286), .ZN(
        u5_mult_82_ab_23__28_) );
  NOR2_X1 u5_mult_82_U2473 ( .A1(u5_mult_82_n386), .A2(u5_mult_82_n286), .ZN(
        u5_mult_82_ab_23__29_) );
  NOR2_X1 u5_mult_82_U2472 ( .A1(u5_mult_82_n442), .A2(u5_mult_82_n286), .ZN(
        u5_mult_82_ab_23__2_) );
  NOR2_X1 u5_mult_82_U2471 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n286), .ZN(
        u5_mult_82_ab_23__30_) );
  NOR2_X1 u5_mult_82_U2470 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n286), .ZN(
        u5_mult_82_ab_23__31_) );
  NOR2_X1 u5_mult_82_U2469 ( .A1(u5_mult_82_n380), .A2(u5_mult_82_n286), .ZN(
        u5_mult_82_ab_23__32_) );
  NOR2_X1 u5_mult_82_U2468 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n286), .ZN(
        u5_mult_82_ab_23__33_) );
  NOR2_X1 u5_mult_82_U2467 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n286), .ZN(
        u5_mult_82_ab_23__34_) );
  NOR2_X1 u5_mult_82_U2466 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n286), .ZN(
        u5_mult_82_ab_23__35_) );
  NOR2_X1 u5_mult_82_U2465 ( .A1(u5_mult_82_n474), .A2(u5_mult_82_n286), .ZN(
        u5_mult_82_ab_23__36_) );
  NOR2_X1 u5_mult_82_U2464 ( .A1(u5_mult_82_n370), .A2(u5_mult_82_n286), .ZN(
        u5_mult_82_ab_23__37_) );
  NOR2_X1 u5_mult_82_U2463 ( .A1(u5_mult_82_n369), .A2(u5_mult_82_n286), .ZN(
        u5_mult_82_ab_23__38_) );
  NOR2_X1 u5_mult_82_U2462 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n286), .ZN(
        u5_mult_82_ab_23__39_) );
  NOR2_X1 u5_mult_82_U2461 ( .A1(u5_mult_82_n440), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__3_) );
  NOR2_X1 u5_mult_82_U2460 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__40_) );
  NOR2_X1 u5_mult_82_U2459 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__41_) );
  NOR2_X1 u5_mult_82_U2458 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__42_) );
  NOR2_X1 u5_mult_82_U2457 ( .A1(u5_mult_82_n356), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__43_) );
  NOR2_X1 u5_mult_82_U2456 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__44_) );
  NOR2_X1 u5_mult_82_U2455 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__45_) );
  NOR2_X1 u5_mult_82_U2454 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__46_) );
  NOR2_X1 u5_mult_82_U2453 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__47_) );
  NOR2_X1 u5_mult_82_U2452 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__48_) );
  NOR2_X1 u5_mult_82_U2451 ( .A1(u5_mult_82_n343), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__49_) );
  NOR2_X1 u5_mult_82_U2450 ( .A1(u5_mult_82_n438), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__4_) );
  NOR2_X1 u5_mult_82_U2449 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__50_) );
  NOR2_X1 u5_mult_82_U2448 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__51_) );
  NOR2_X1 u5_mult_82_U2447 ( .A1(u5_mult_82_n336), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__52_) );
  NOR2_X1 u5_mult_82_U2446 ( .A1(u5_mult_82_n436), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__5_) );
  NOR2_X1 u5_mult_82_U2445 ( .A1(u5_mult_82_n434), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__6_) );
  NOR2_X1 u5_mult_82_U2444 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__7_) );
  NOR2_X1 u5_mult_82_U2443 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__8_) );
  NOR2_X1 u5_mult_82_U2442 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n287), .ZN(
        u5_mult_82_ab_23__9_) );
  NOR2_X1 u5_mult_82_U2441 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__0_) );
  NOR2_X1 u5_mult_82_U2440 ( .A1(u5_mult_82_n477), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__10_) );
  NOR2_X1 u5_mult_82_U2439 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__11_) );
  NOR2_X1 u5_mult_82_U2438 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__12_) );
  NOR2_X1 u5_mult_82_U2437 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__13_) );
  NOR2_X1 u5_mult_82_U2436 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__14_) );
  NOR2_X1 u5_mult_82_U2435 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__15_) );
  NOR2_X1 u5_mult_82_U2434 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__16_) );
  NOR2_X1 u5_mult_82_U2433 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__17_) );
  NOR2_X1 u5_mult_82_U2432 ( .A1(u5_mult_82_n406), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__18_) );
  NOR2_X1 u5_mult_82_U2431 ( .A1(u5_mult_82_n404), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__19_) );
  NOR2_X1 u5_mult_82_U2430 ( .A1(u5_mult_82_n443), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__1_) );
  NOR2_X1 u5_mult_82_U2429 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__20_) );
  NOR2_X1 u5_mult_82_U2428 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__21_) );
  NOR2_X1 u5_mult_82_U2427 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__22_) );
  NOR2_X1 u5_mult_82_U2426 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__23_) );
  NOR2_X1 u5_mult_82_U2425 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n284), .ZN(
        u5_mult_82_ab_24__24_) );
  NOR2_X1 u5_mult_82_U2424 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n284), .ZN(
        u5_mult_82_ab_24__25_) );
  NOR2_X1 u5_mult_82_U2423 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n284), .ZN(
        u5_mult_82_ab_24__26_) );
  NOR2_X1 u5_mult_82_U2422 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n284), .ZN(
        u5_mult_82_ab_24__27_) );
  NOR2_X1 u5_mult_82_U2421 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n284), .ZN(
        u5_mult_82_ab_24__28_) );
  NOR2_X1 u5_mult_82_U2420 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n284), .ZN(
        u5_mult_82_ab_24__29_) );
  NOR2_X1 u5_mult_82_U2419 ( .A1(u5_mult_82_n442), .A2(u5_mult_82_n284), .ZN(
        u5_mult_82_ab_24__2_) );
  NOR2_X1 u5_mult_82_U2418 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n284), .ZN(
        u5_mult_82_ab_24__30_) );
  NOR2_X1 u5_mult_82_U2417 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n284), .ZN(
        u5_mult_82_ab_24__31_) );
  NOR2_X1 u5_mult_82_U2416 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n284), .ZN(
        u5_mult_82_ab_24__32_) );
  NOR2_X1 u5_mult_82_U2415 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n284), .ZN(
        u5_mult_82_ab_24__33_) );
  NOR2_X1 u5_mult_82_U2414 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n284), .ZN(
        u5_mult_82_ab_24__34_) );
  NOR2_X1 u5_mult_82_U2413 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n284), .ZN(
        u5_mult_82_ab_24__35_) );
  NOR2_X1 u5_mult_82_U2412 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n284), .ZN(
        u5_mult_82_ab_24__36_) );
  NOR2_X1 u5_mult_82_U2411 ( .A1(u5_mult_82_n370), .A2(u5_mult_82_n284), .ZN(
        u5_mult_82_ab_24__37_) );
  NOR2_X1 u5_mult_82_U2410 ( .A1(u5_mult_82_n369), .A2(u5_mult_82_n284), .ZN(
        u5_mult_82_ab_24__38_) );
  NOR2_X1 u5_mult_82_U2409 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n284), .ZN(
        u5_mult_82_ab_24__39_) );
  NOR2_X1 u5_mult_82_U2408 ( .A1(u5_mult_82_n440), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__3_) );
  NOR2_X1 u5_mult_82_U2407 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__40_) );
  NOR2_X1 u5_mult_82_U2406 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__41_) );
  NOR2_X1 u5_mult_82_U2405 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__42_) );
  NOR2_X1 u5_mult_82_U2404 ( .A1(u5_mult_82_n356), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__43_) );
  NOR2_X1 u5_mult_82_U2403 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__44_) );
  NOR2_X1 u5_mult_82_U2402 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__45_) );
  NOR2_X1 u5_mult_82_U2401 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__46_) );
  NOR2_X1 u5_mult_82_U2400 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__47_) );
  NOR2_X1 u5_mult_82_U2399 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__48_) );
  NOR2_X1 u5_mult_82_U2398 ( .A1(u5_mult_82_n343), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__49_) );
  NOR2_X1 u5_mult_82_U2397 ( .A1(u5_mult_82_n438), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__4_) );
  NOR2_X1 u5_mult_82_U2396 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__50_) );
  NOR2_X1 u5_mult_82_U2395 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__51_) );
  NOR2_X1 u5_mult_82_U2394 ( .A1(u5_mult_82_n336), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__52_) );
  NOR2_X1 u5_mult_82_U2393 ( .A1(u5_mult_82_n436), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__5_) );
  NOR2_X1 u5_mult_82_U2392 ( .A1(u5_mult_82_n434), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__6_) );
  NOR2_X1 u5_mult_82_U2391 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__7_) );
  NOR2_X1 u5_mult_82_U2390 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__8_) );
  NOR2_X1 u5_mult_82_U2389 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n285), .ZN(
        u5_mult_82_ab_24__9_) );
  NOR2_X1 u5_mult_82_U2388 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__0_) );
  NOR2_X1 u5_mult_82_U2387 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__10_) );
  NOR2_X1 u5_mult_82_U2386 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__11_) );
  NOR2_X1 u5_mult_82_U2385 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__12_) );
  NOR2_X1 u5_mult_82_U2384 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__13_) );
  NOR2_X1 u5_mult_82_U2383 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__14_) );
  NOR2_X1 u5_mult_82_U2382 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__15_) );
  NOR2_X1 u5_mult_82_U2381 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__16_) );
  NOR2_X1 u5_mult_82_U2380 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__17_) );
  NOR2_X1 u5_mult_82_U2379 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__18_) );
  NOR2_X1 u5_mult_82_U2378 ( .A1(u5_mult_82_n404), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__19_) );
  NOR2_X1 u5_mult_82_U2377 ( .A1(u5_mult_82_n443), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__1_) );
  NOR2_X1 u5_mult_82_U2376 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__20_) );
  NOR2_X1 u5_mult_82_U2375 ( .A1(u5_mult_82_n402), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__21_) );
  NOR2_X1 u5_mult_82_U2374 ( .A1(u5_mult_82_n400), .A2(u5_mult_82_n462), .ZN(
        u5_mult_82_ab_25__22_) );
  NOR2_X1 u5_mult_82_U2373 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n462), .ZN(
        u5_mult_82_ab_25__23_) );
  NOR2_X1 u5_mult_82_U2372 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n462), .ZN(
        u5_mult_82_ab_25__24_) );
  NOR2_X1 u5_mult_82_U2371 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n462), .ZN(
        u5_mult_82_ab_25__25_) );
  NOR2_X1 u5_mult_82_U2370 ( .A1(u5_mult_82_n392), .A2(u5_mult_82_n282), .ZN(
        u5_mult_82_ab_25__26_) );
  NOR2_X1 u5_mult_82_U2369 ( .A1(u5_mult_82_n390), .A2(u5_mult_82_n282), .ZN(
        u5_mult_82_ab_25__27_) );
  NOR2_X1 u5_mult_82_U2368 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n462), .ZN(
        u5_mult_82_ab_25__28_) );
  NOR2_X1 u5_mult_82_U2367 ( .A1(u5_mult_82_n386), .A2(u5_mult_82_n462), .ZN(
        u5_mult_82_ab_25__29_) );
  NOR2_X1 u5_mult_82_U2366 ( .A1(u5_mult_82_n442), .A2(u5_mult_82_n282), .ZN(
        u5_mult_82_ab_25__2_) );
  NOR2_X1 u5_mult_82_U2365 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n282), .ZN(
        u5_mult_82_ab_25__30_) );
  NOR2_X1 u5_mult_82_U2364 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n282), .ZN(
        u5_mult_82_ab_25__31_) );
  NOR2_X1 u5_mult_82_U2363 ( .A1(u5_mult_82_n380), .A2(u5_mult_82_n282), .ZN(
        u5_mult_82_ab_25__32_) );
  NOR2_X1 u5_mult_82_U2362 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n282), .ZN(
        u5_mult_82_ab_25__33_) );
  NOR2_X1 u5_mult_82_U2361 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n282), .ZN(
        u5_mult_82_ab_25__34_) );
  NOR2_X1 u5_mult_82_U2360 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n282), .ZN(
        u5_mult_82_ab_25__35_) );
  NOR2_X1 u5_mult_82_U2359 ( .A1(u5_mult_82_n474), .A2(u5_mult_82_n282), .ZN(
        u5_mult_82_ab_25__36_) );
  NOR2_X1 u5_mult_82_U2358 ( .A1(u5_mult_82_n370), .A2(u5_mult_82_n282), .ZN(
        u5_mult_82_ab_25__37_) );
  NOR2_X1 u5_mult_82_U2357 ( .A1(u5_mult_82_n369), .A2(u5_mult_82_n282), .ZN(
        u5_mult_82_ab_25__38_) );
  NOR2_X1 u5_mult_82_U2356 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n282), .ZN(
        u5_mult_82_ab_25__39_) );
  NOR2_X1 u5_mult_82_U2355 ( .A1(u5_mult_82_n440), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__3_) );
  NOR2_X1 u5_mult_82_U2354 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__40_) );
  NOR2_X1 u5_mult_82_U2353 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__41_) );
  NOR2_X1 u5_mult_82_U2352 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__42_) );
  NOR2_X1 u5_mult_82_U2351 ( .A1(u5_mult_82_n356), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__43_) );
  NOR2_X1 u5_mult_82_U2350 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__44_) );
  NOR2_X1 u5_mult_82_U2349 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__45_) );
  NOR2_X1 u5_mult_82_U2348 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__46_) );
  NOR2_X1 u5_mult_82_U2347 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__47_) );
  NOR2_X1 u5_mult_82_U2346 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__48_) );
  NOR2_X1 u5_mult_82_U2345 ( .A1(u5_mult_82_n343), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__49_) );
  NOR2_X1 u5_mult_82_U2344 ( .A1(u5_mult_82_n438), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__4_) );
  NOR2_X1 u5_mult_82_U2343 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__50_) );
  NOR2_X1 u5_mult_82_U2342 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__51_) );
  NOR2_X1 u5_mult_82_U2341 ( .A1(u5_mult_82_n336), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__52_) );
  NOR2_X1 u5_mult_82_U2340 ( .A1(u5_mult_82_n436), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__5_) );
  NOR2_X1 u5_mult_82_U2339 ( .A1(u5_mult_82_n434), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__6_) );
  NOR2_X1 u5_mult_82_U2338 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__7_) );
  NOR2_X1 u5_mult_82_U2337 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__8_) );
  NOR2_X1 u5_mult_82_U2336 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n283), .ZN(
        u5_mult_82_ab_25__9_) );
  NOR2_X1 u5_mult_82_U2335 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__0_) );
  NOR2_X1 u5_mult_82_U2334 ( .A1(u5_mult_82_n477), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__10_) );
  NOR2_X1 u5_mult_82_U2333 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__11_) );
  NOR2_X1 u5_mult_82_U2332 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__12_) );
  NOR2_X1 u5_mult_82_U2331 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__13_) );
  NOR2_X1 u5_mult_82_U2330 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__14_) );
  NOR2_X1 u5_mult_82_U2329 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__15_) );
  NOR2_X1 u5_mult_82_U2328 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__16_) );
  NOR2_X1 u5_mult_82_U2327 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__17_) );
  NOR2_X1 u5_mult_82_U2326 ( .A1(u5_mult_82_n476), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__18_) );
  NOR2_X1 u5_mult_82_U2325 ( .A1(u5_mult_82_n404), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__19_) );
  NOR2_X1 u5_mult_82_U2324 ( .A1(u5_mult_82_n443), .A2(u5_mult_82_n281), .ZN(
        u5_mult_82_ab_26__1_) );
  NOR2_X1 u5_mult_82_U2323 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n281), .ZN(
        u5_mult_82_ab_26__20_) );
  NOR2_X1 u5_mult_82_U2322 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n281), .ZN(
        u5_mult_82_ab_26__21_) );
  NOR2_X1 u5_mult_82_U2321 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n281), .ZN(
        u5_mult_82_ab_26__22_) );
  NOR2_X1 u5_mult_82_U2320 ( .A1(u5_mult_82_n398), .A2(u5_mult_82_n281), .ZN(
        u5_mult_82_ab_26__23_) );
  NOR2_X1 u5_mult_82_U2319 ( .A1(u5_mult_82_n396), .A2(u5_mult_82_n281), .ZN(
        u5_mult_82_ab_26__24_) );
  NOR2_X1 u5_mult_82_U2318 ( .A1(u5_mult_82_n394), .A2(u5_mult_82_n281), .ZN(
        u5_mult_82_ab_26__25_) );
  NOR2_X1 u5_mult_82_U2317 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n281), .ZN(
        u5_mult_82_ab_26__26_) );
  NOR2_X1 u5_mult_82_U2316 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n281), .ZN(
        u5_mult_82_ab_26__27_) );
  NOR2_X1 u5_mult_82_U2315 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n281), .ZN(
        u5_mult_82_ab_26__28_) );
  NOR2_X1 u5_mult_82_U2314 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n281), .ZN(
        u5_mult_82_ab_26__29_) );
  NOR2_X1 u5_mult_82_U2313 ( .A1(u5_mult_82_n442), .A2(u5_mult_82_n281), .ZN(
        u5_mult_82_ab_26__2_) );
  NOR2_X1 u5_mult_82_U2312 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n281), .ZN(
        u5_mult_82_ab_26__30_) );
  NOR2_X1 u5_mult_82_U2311 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n281), .ZN(
        u5_mult_82_ab_26__31_) );
  NOR2_X1 u5_mult_82_U2310 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n281), .ZN(
        u5_mult_82_ab_26__32_) );
  NOR2_X1 u5_mult_82_U2309 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n281), .ZN(
        u5_mult_82_ab_26__33_) );
  NOR2_X1 u5_mult_82_U2308 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n281), .ZN(
        u5_mult_82_ab_26__34_) );
  NOR2_X1 u5_mult_82_U2307 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n281), .ZN(
        u5_mult_82_ab_26__35_) );
  NOR2_X1 u5_mult_82_U2306 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n281), .ZN(
        u5_mult_82_ab_26__36_) );
  NOR2_X1 u5_mult_82_U2305 ( .A1(u5_mult_82_n370), .A2(u5_mult_82_n281), .ZN(
        u5_mult_82_ab_26__37_) );
  NOR2_X1 u5_mult_82_U2304 ( .A1(u5_mult_82_n369), .A2(u5_mult_82_n281), .ZN(
        u5_mult_82_ab_26__38_) );
  NOR2_X1 u5_mult_82_U2303 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n281), .ZN(
        u5_mult_82_ab_26__39_) );
  NOR2_X1 u5_mult_82_U2302 ( .A1(u5_mult_82_n440), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__3_) );
  NOR2_X1 u5_mult_82_U2301 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__40_) );
  NOR2_X1 u5_mult_82_U2300 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__41_) );
  NOR2_X1 u5_mult_82_U2299 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__42_) );
  NOR2_X1 u5_mult_82_U2298 ( .A1(u5_mult_82_n356), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__43_) );
  NOR2_X1 u5_mult_82_U2297 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__44_) );
  NOR2_X1 u5_mult_82_U2296 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__45_) );
  NOR2_X1 u5_mult_82_U2295 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__46_) );
  NOR2_X1 u5_mult_82_U2294 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__47_) );
  NOR2_X1 u5_mult_82_U2293 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__48_) );
  NOR2_X1 u5_mult_82_U2292 ( .A1(u5_mult_82_n343), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__49_) );
  NOR2_X1 u5_mult_82_U2291 ( .A1(u5_mult_82_n438), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__4_) );
  NOR2_X1 u5_mult_82_U2290 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__50_) );
  NOR2_X1 u5_mult_82_U2289 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__51_) );
  NOR2_X1 u5_mult_82_U2288 ( .A1(u5_mult_82_n336), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__52_) );
  NOR2_X1 u5_mult_82_U2287 ( .A1(u5_mult_82_n436), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__5_) );
  NOR2_X1 u5_mult_82_U2286 ( .A1(u5_mult_82_n434), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__6_) );
  NOR2_X1 u5_mult_82_U2285 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__7_) );
  NOR2_X1 u5_mult_82_U2284 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__8_) );
  NOR2_X1 u5_mult_82_U2283 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n280), .ZN(
        u5_mult_82_ab_26__9_) );
  NOR2_X1 u5_mult_82_U2282 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n279), .ZN(
        u5_mult_82_ab_27__0_) );
  NOR2_X1 u5_mult_82_U2281 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n278), .ZN(
        u5_mult_82_ab_27__10_) );
  NOR2_X1 u5_mult_82_U2280 ( .A1(u5_mult_82_n426), .A2(u5_mult_82_n278), .ZN(
        u5_mult_82_ab_27__11_) );
  NOR2_X1 u5_mult_82_U2279 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n278), .ZN(
        u5_mult_82_ab_27__12_) );
  NOR2_X1 u5_mult_82_U2278 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n278), .ZN(
        u5_mult_82_ab_27__13_) );
  NOR2_X1 u5_mult_82_U2277 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n278), .ZN(
        u5_mult_82_ab_27__14_) );
  NOR2_X1 u5_mult_82_U2276 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n279), .ZN(
        u5_mult_82_ab_27__15_) );
  NOR2_X1 u5_mult_82_U2275 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n279), .ZN(
        u5_mult_82_ab_27__16_) );
  NOR2_X1 u5_mult_82_U2274 ( .A1(u5_mult_82_n409), .A2(u5_mult_82_n278), .ZN(
        u5_mult_82_ab_27__17_) );
  NOR2_X1 u5_mult_82_U2273 ( .A1(u5_mult_82_n476), .A2(u5_mult_82_n278), .ZN(
        u5_mult_82_ab_27__18_) );
  NOR2_X1 u5_mult_82_U2272 ( .A1(u5_mult_82_n404), .A2(u5_mult_82_n278), .ZN(
        u5_mult_82_ab_27__19_) );
  NOR2_X1 u5_mult_82_U2271 ( .A1(u5_mult_82_n443), .A2(u5_mult_82_n279), .ZN(
        u5_mult_82_ab_27__1_) );
  NOR2_X1 u5_mult_82_U2270 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n278), .ZN(
        u5_mult_82_ab_27__20_) );
  NOR2_X1 u5_mult_82_U2269 ( .A1(u5_mult_82_n402), .A2(u5_mult_82_n461), .ZN(
        u5_mult_82_ab_27__21_) );
  NOR2_X1 u5_mult_82_U2268 ( .A1(u5_mult_82_n400), .A2(u5_mult_82_n461), .ZN(
        u5_mult_82_ab_27__22_) );
  NOR2_X1 u5_mult_82_U2267 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n461), .ZN(
        u5_mult_82_ab_27__23_) );
  NOR2_X1 u5_mult_82_U2266 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n461), .ZN(
        u5_mult_82_ab_27__24_) );
  NOR2_X1 u5_mult_82_U2265 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n461), .ZN(
        u5_mult_82_ab_27__25_) );
  NOR2_X1 u5_mult_82_U2264 ( .A1(u5_mult_82_n392), .A2(u5_mult_82_n461), .ZN(
        u5_mult_82_ab_27__26_) );
  NOR2_X1 u5_mult_82_U2263 ( .A1(u5_mult_82_n390), .A2(u5_mult_82_n461), .ZN(
        u5_mult_82_ab_27__27_) );
  NOR2_X1 u5_mult_82_U2262 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n461), .ZN(
        u5_mult_82_ab_27__28_) );
  NOR2_X1 u5_mult_82_U2261 ( .A1(u5_mult_82_n386), .A2(u5_mult_82_n461), .ZN(
        u5_mult_82_ab_27__29_) );
  NOR2_X1 u5_mult_82_U2260 ( .A1(u5_mult_82_n442), .A2(u5_mult_82_n278), .ZN(
        u5_mult_82_ab_27__2_) );
  NOR2_X1 u5_mult_82_U2259 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n278), .ZN(
        u5_mult_82_ab_27__30_) );
  NOR2_X1 u5_mult_82_U2258 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n278), .ZN(
        u5_mult_82_ab_27__31_) );
  NOR2_X1 u5_mult_82_U2257 ( .A1(u5_mult_82_n380), .A2(u5_mult_82_n278), .ZN(
        u5_mult_82_ab_27__32_) );
  NOR2_X1 u5_mult_82_U2256 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n278), .ZN(
        u5_mult_82_ab_27__33_) );
  NOR2_X1 u5_mult_82_U2255 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n278), .ZN(
        u5_mult_82_ab_27__34_) );
  NOR2_X1 u5_mult_82_U2254 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n278), .ZN(
        u5_mult_82_ab_27__35_) );
  NOR2_X1 u5_mult_82_U2253 ( .A1(u5_mult_82_n474), .A2(u5_mult_82_n278), .ZN(
        u5_mult_82_ab_27__36_) );
  NOR2_X1 u5_mult_82_U2252 ( .A1(u5_mult_82_n370), .A2(u5_mult_82_n278), .ZN(
        u5_mult_82_ab_27__37_) );
  NOR2_X1 u5_mult_82_U2251 ( .A1(u5_mult_82_n369), .A2(u5_mult_82_n278), .ZN(
        u5_mult_82_ab_27__38_) );
  NOR2_X1 u5_mult_82_U2250 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n278), .ZN(
        u5_mult_82_ab_27__39_) );
  NOR2_X1 u5_mult_82_U2249 ( .A1(u5_mult_82_n440), .A2(u5_mult_82_n279), .ZN(
        u5_mult_82_ab_27__3_) );
  NOR2_X1 u5_mult_82_U2248 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n279), .ZN(
        u5_mult_82_ab_27__40_) );
  NOR2_X1 u5_mult_82_U2247 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n279), .ZN(
        u5_mult_82_ab_27__41_) );
  NOR2_X1 u5_mult_82_U2246 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n279), .ZN(
        u5_mult_82_ab_27__42_) );
  NOR2_X1 u5_mult_82_U2245 ( .A1(u5_mult_82_n356), .A2(u5_mult_82_n279), .ZN(
        u5_mult_82_ab_27__43_) );
  NOR2_X1 u5_mult_82_U2244 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n279), .ZN(
        u5_mult_82_ab_27__44_) );
  NOR2_X1 u5_mult_82_U2243 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n279), .ZN(
        u5_mult_82_ab_27__45_) );
  NOR2_X1 u5_mult_82_U2242 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n279), .ZN(
        u5_mult_82_ab_27__46_) );
  NOR2_X1 u5_mult_82_U2241 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n279), .ZN(
        u5_mult_82_ab_27__47_) );
  NOR2_X1 u5_mult_82_U2240 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n279), .ZN(
        u5_mult_82_ab_27__48_) );
  NOR2_X1 u5_mult_82_U2239 ( .A1(u5_mult_82_n343), .A2(u5_mult_82_n279), .ZN(
        u5_mult_82_ab_27__49_) );
  NOR2_X1 u5_mult_82_U2238 ( .A1(u5_mult_82_n438), .A2(u5_mult_82_n279), .ZN(
        u5_mult_82_ab_27__4_) );
  NOR2_X1 u5_mult_82_U2237 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n279), .ZN(
        u5_mult_82_ab_27__50_) );
  NOR2_X1 u5_mult_82_U2236 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n279), .ZN(
        u5_mult_82_ab_27__51_) );
  NOR2_X1 u5_mult_82_U2235 ( .A1(u5_mult_82_n336), .A2(u5_mult_82_n279), .ZN(
        u5_mult_82_ab_27__52_) );
  NOR2_X1 u5_mult_82_U2234 ( .A1(u5_mult_82_n436), .A2(u5_mult_82_n279), .ZN(
        u5_mult_82_ab_27__5_) );
  NOR2_X1 u5_mult_82_U2233 ( .A1(u5_mult_82_n434), .A2(u5_mult_82_n279), .ZN(
        u5_mult_82_ab_27__6_) );
  NOR2_X1 u5_mult_82_U2232 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n279), .ZN(
        u5_mult_82_ab_27__7_) );
  NOR2_X1 u5_mult_82_U2231 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n279), .ZN(
        u5_mult_82_ab_27__8_) );
  NOR2_X1 u5_mult_82_U2230 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n279), .ZN(
        u5_mult_82_ab_27__9_) );
  NOR2_X1 u5_mult_82_U2229 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n276), .ZN(
        u5_mult_82_ab_28__0_) );
  NOR2_X1 u5_mult_82_U2228 ( .A1(u5_mult_82_n477), .A2(u5_mult_82_n275), .ZN(
        u5_mult_82_ab_28__10_) );
  NOR2_X1 u5_mult_82_U2227 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n275), .ZN(
        u5_mult_82_ab_28__11_) );
  NOR2_X1 u5_mult_82_U2226 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n275), .ZN(
        u5_mult_82_ab_28__12_) );
  NOR2_X1 u5_mult_82_U2225 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n275), .ZN(
        u5_mult_82_ab_28__13_) );
  NOR2_X1 u5_mult_82_U2224 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n275), .ZN(
        u5_mult_82_ab_28__14_) );
  NOR2_X1 u5_mult_82_U2223 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n276), .ZN(
        u5_mult_82_ab_28__15_) );
  NOR2_X1 u5_mult_82_U2222 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n276), .ZN(
        u5_mult_82_ab_28__16_) );
  NOR2_X1 u5_mult_82_U2221 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n275), .ZN(
        u5_mult_82_ab_28__17_) );
  NOR2_X1 u5_mult_82_U2220 ( .A1(u5_mult_82_n476), .A2(u5_mult_82_n275), .ZN(
        u5_mult_82_ab_28__18_) );
  NOR2_X1 u5_mult_82_U2219 ( .A1(u5_mult_82_n404), .A2(u5_mult_82_n275), .ZN(
        u5_mult_82_ab_28__19_) );
  NOR2_X1 u5_mult_82_U2218 ( .A1(u5_mult_82_n443), .A2(u5_mult_82_n276), .ZN(
        u5_mult_82_ab_28__1_) );
  NOR2_X1 u5_mult_82_U2217 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n276), .ZN(
        u5_mult_82_ab_28__20_) );
  NOR2_X1 u5_mult_82_U2216 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n275), .ZN(
        u5_mult_82_ab_28__21_) );
  NOR2_X1 u5_mult_82_U2215 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n277), .ZN(
        u5_mult_82_ab_28__22_) );
  NOR2_X1 u5_mult_82_U2214 ( .A1(u5_mult_82_n398), .A2(u5_mult_82_n277), .ZN(
        u5_mult_82_ab_28__23_) );
  NOR2_X1 u5_mult_82_U2213 ( .A1(u5_mult_82_n396), .A2(u5_mult_82_n277), .ZN(
        u5_mult_82_ab_28__24_) );
  NOR2_X1 u5_mult_82_U2212 ( .A1(u5_mult_82_n394), .A2(u5_mult_82_n277), .ZN(
        u5_mult_82_ab_28__25_) );
  NOR2_X1 u5_mult_82_U2211 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n277), .ZN(
        u5_mult_82_ab_28__26_) );
  NOR2_X1 u5_mult_82_U2210 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n277), .ZN(
        u5_mult_82_ab_28__27_) );
  NOR2_X1 u5_mult_82_U2209 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n277), .ZN(
        u5_mult_82_ab_28__28_) );
  NOR2_X1 u5_mult_82_U2208 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n275), .ZN(
        u5_mult_82_ab_28__29_) );
  NOR2_X1 u5_mult_82_U2207 ( .A1(u5_mult_82_n442), .A2(u5_mult_82_n275), .ZN(
        u5_mult_82_ab_28__2_) );
  NOR2_X1 u5_mult_82_U2206 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n275), .ZN(
        u5_mult_82_ab_28__30_) );
  NOR2_X1 u5_mult_82_U2205 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n275), .ZN(
        u5_mult_82_ab_28__31_) );
  NOR2_X1 u5_mult_82_U2204 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n275), .ZN(
        u5_mult_82_ab_28__32_) );
  NOR2_X1 u5_mult_82_U2203 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n275), .ZN(
        u5_mult_82_ab_28__33_) );
  NOR2_X1 u5_mult_82_U2202 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n275), .ZN(
        u5_mult_82_ab_28__34_) );
  NOR2_X1 u5_mult_82_U2201 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n275), .ZN(
        u5_mult_82_ab_28__35_) );
  NOR2_X1 u5_mult_82_U2200 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n275), .ZN(
        u5_mult_82_ab_28__36_) );
  NOR2_X1 u5_mult_82_U2199 ( .A1(u5_mult_82_n370), .A2(u5_mult_82_n275), .ZN(
        u5_mult_82_ab_28__37_) );
  NOR2_X1 u5_mult_82_U2198 ( .A1(u5_mult_82_n369), .A2(u5_mult_82_n275), .ZN(
        u5_mult_82_ab_28__38_) );
  NOR2_X1 u5_mult_82_U2197 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n275), .ZN(
        u5_mult_82_ab_28__39_) );
  NOR2_X1 u5_mult_82_U2196 ( .A1(u5_mult_82_n440), .A2(u5_mult_82_n276), .ZN(
        u5_mult_82_ab_28__3_) );
  NOR2_X1 u5_mult_82_U2195 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n276), .ZN(
        u5_mult_82_ab_28__40_) );
  NOR2_X1 u5_mult_82_U2194 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n276), .ZN(
        u5_mult_82_ab_28__41_) );
  NOR2_X1 u5_mult_82_U2193 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n276), .ZN(
        u5_mult_82_ab_28__42_) );
  NOR2_X1 u5_mult_82_U2192 ( .A1(u5_mult_82_n356), .A2(u5_mult_82_n276), .ZN(
        u5_mult_82_ab_28__43_) );
  NOR2_X1 u5_mult_82_U2191 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n276), .ZN(
        u5_mult_82_ab_28__44_) );
  NOR2_X1 u5_mult_82_U2190 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n276), .ZN(
        u5_mult_82_ab_28__45_) );
  NOR2_X1 u5_mult_82_U2189 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n276), .ZN(
        u5_mult_82_ab_28__46_) );
  NOR2_X1 u5_mult_82_U2188 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n276), .ZN(
        u5_mult_82_ab_28__47_) );
  NOR2_X1 u5_mult_82_U2187 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n276), .ZN(
        u5_mult_82_ab_28__48_) );
  NOR2_X1 u5_mult_82_U2186 ( .A1(u5_mult_82_n343), .A2(u5_mult_82_n276), .ZN(
        u5_mult_82_ab_28__49_) );
  NOR2_X1 u5_mult_82_U2185 ( .A1(u5_mult_82_n438), .A2(u5_mult_82_n276), .ZN(
        u5_mult_82_ab_28__4_) );
  NOR2_X1 u5_mult_82_U2184 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n276), .ZN(
        u5_mult_82_ab_28__50_) );
  NOR2_X1 u5_mult_82_U2183 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n276), .ZN(
        u5_mult_82_ab_28__51_) );
  NOR2_X1 u5_mult_82_U2182 ( .A1(u5_mult_82_n336), .A2(u5_mult_82_n276), .ZN(
        u5_mult_82_ab_28__52_) );
  NOR2_X1 u5_mult_82_U2181 ( .A1(u5_mult_82_n436), .A2(u5_mult_82_n276), .ZN(
        u5_mult_82_ab_28__5_) );
  NOR2_X1 u5_mult_82_U2180 ( .A1(u5_mult_82_n434), .A2(u5_mult_82_n276), .ZN(
        u5_mult_82_ab_28__6_) );
  NOR2_X1 u5_mult_82_U2179 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n276), .ZN(
        u5_mult_82_ab_28__7_) );
  NOR2_X1 u5_mult_82_U2178 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n276), .ZN(
        u5_mult_82_ab_28__8_) );
  NOR2_X1 u5_mult_82_U2177 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n276), .ZN(
        u5_mult_82_ab_28__9_) );
  NOR2_X1 u5_mult_82_U2176 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__0_) );
  NOR2_X1 u5_mult_82_U2175 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n272), .ZN(
        u5_mult_82_ab_29__10_) );
  NOR2_X1 u5_mult_82_U2174 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__11_) );
  NOR2_X1 u5_mult_82_U2173 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n272), .ZN(
        u5_mult_82_ab_29__12_) );
  NOR2_X1 u5_mult_82_U2172 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__13_) );
  NOR2_X1 u5_mult_82_U2171 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__14_) );
  NOR2_X1 u5_mult_82_U2170 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__15_) );
  NOR2_X1 u5_mult_82_U2169 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__16_) );
  NOR2_X1 u5_mult_82_U2168 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__17_) );
  NOR2_X1 u5_mult_82_U2167 ( .A1(u5_mult_82_n476), .A2(u5_mult_82_n272), .ZN(
        u5_mult_82_ab_29__18_) );
  NOR2_X1 u5_mult_82_U2166 ( .A1(u5_mult_82_n404), .A2(u5_mult_82_n272), .ZN(
        u5_mult_82_ab_29__19_) );
  NOR2_X1 u5_mult_82_U2165 ( .A1(u5_mult_82_n443), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__1_) );
  NOR2_X1 u5_mult_82_U2164 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n272), .ZN(
        u5_mult_82_ab_29__20_) );
  NOR2_X1 u5_mult_82_U2163 ( .A1(u5_mult_82_n402), .A2(u5_mult_82_n274), .ZN(
        u5_mult_82_ab_29__21_) );
  NOR2_X1 u5_mult_82_U2162 ( .A1(u5_mult_82_n400), .A2(u5_mult_82_n274), .ZN(
        u5_mult_82_ab_29__22_) );
  NOR2_X1 u5_mult_82_U2161 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n274), .ZN(
        u5_mult_82_ab_29__23_) );
  NOR2_X1 u5_mult_82_U2160 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n274), .ZN(
        u5_mult_82_ab_29__24_) );
  NOR2_X1 u5_mult_82_U2159 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n274), .ZN(
        u5_mult_82_ab_29__25_) );
  NOR2_X1 u5_mult_82_U2158 ( .A1(u5_mult_82_n392), .A2(u5_mult_82_n274), .ZN(
        u5_mult_82_ab_29__26_) );
  NOR2_X1 u5_mult_82_U2157 ( .A1(u5_mult_82_n390), .A2(u5_mult_82_n272), .ZN(
        u5_mult_82_ab_29__27_) );
  NOR2_X1 u5_mult_82_U2156 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__28_) );
  NOR2_X1 u5_mult_82_U2155 ( .A1(u5_mult_82_n386), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__29_) );
  NOR2_X1 u5_mult_82_U2154 ( .A1(u5_mult_82_n442), .A2(u5_mult_82_n272), .ZN(
        u5_mult_82_ab_29__2_) );
  NOR2_X1 u5_mult_82_U2153 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n272), .ZN(
        u5_mult_82_ab_29__30_) );
  NOR2_X1 u5_mult_82_U2152 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n272), .ZN(
        u5_mult_82_ab_29__31_) );
  NOR2_X1 u5_mult_82_U2151 ( .A1(u5_mult_82_n380), .A2(u5_mult_82_n272), .ZN(
        u5_mult_82_ab_29__32_) );
  NOR2_X1 u5_mult_82_U2150 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n272), .ZN(
        u5_mult_82_ab_29__33_) );
  NOR2_X1 u5_mult_82_U2149 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n272), .ZN(
        u5_mult_82_ab_29__34_) );
  NOR2_X1 u5_mult_82_U2148 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n272), .ZN(
        u5_mult_82_ab_29__35_) );
  NOR2_X1 u5_mult_82_U2147 ( .A1(u5_mult_82_n474), .A2(u5_mult_82_n272), .ZN(
        u5_mult_82_ab_29__36_) );
  NOR2_X1 u5_mult_82_U2146 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n272), .ZN(
        u5_mult_82_ab_29__37_) );
  NOR2_X1 u5_mult_82_U2145 ( .A1(u5_mult_82_n369), .A2(u5_mult_82_n272), .ZN(
        u5_mult_82_ab_29__38_) );
  NOR2_X1 u5_mult_82_U2144 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n272), .ZN(
        u5_mult_82_ab_29__39_) );
  NOR2_X1 u5_mult_82_U2143 ( .A1(u5_mult_82_n440), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__3_) );
  NOR2_X1 u5_mult_82_U2142 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__40_) );
  NOR2_X1 u5_mult_82_U2141 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__41_) );
  NOR2_X1 u5_mult_82_U2140 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__42_) );
  NOR2_X1 u5_mult_82_U2139 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__43_) );
  NOR2_X1 u5_mult_82_U2138 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__44_) );
  NOR2_X1 u5_mult_82_U2137 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__45_) );
  NOR2_X1 u5_mult_82_U2136 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__46_) );
  NOR2_X1 u5_mult_82_U2135 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__47_) );
  NOR2_X1 u5_mult_82_U2134 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__48_) );
  NOR2_X1 u5_mult_82_U2133 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__49_) );
  NOR2_X1 u5_mult_82_U2132 ( .A1(u5_mult_82_n438), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__4_) );
  NOR2_X1 u5_mult_82_U2131 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__50_) );
  NOR2_X1 u5_mult_82_U2130 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__51_) );
  NOR2_X1 u5_mult_82_U2129 ( .A1(u5_mult_82_n336), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__52_) );
  NOR2_X1 u5_mult_82_U2128 ( .A1(u5_mult_82_n436), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__5_) );
  NOR2_X1 u5_mult_82_U2127 ( .A1(u5_mult_82_n434), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__6_) );
  NOR2_X1 u5_mult_82_U2126 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__7_) );
  NOR2_X1 u5_mult_82_U2125 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n273), .ZN(
        u5_mult_82_ab_29__8_) );
  NOR2_X1 u5_mult_82_U2124 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n272), .ZN(
        u5_mult_82_ab_29__9_) );
  NOR2_X1 u5_mult_82_U2123 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__0_) );
  NOR2_X1 u5_mult_82_U2122 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__10_) );
  NOR2_X1 u5_mult_82_U2121 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__11_) );
  NOR2_X1 u5_mult_82_U2120 ( .A1(u5_mult_82_n422), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__12_) );
  NOR2_X1 u5_mult_82_U2119 ( .A1(u5_mult_82_n419), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__13_) );
  NOR2_X1 u5_mult_82_U2118 ( .A1(u5_mult_82_n416), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__14_) );
  NOR2_X1 u5_mult_82_U2117 ( .A1(u5_mult_82_n413), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__15_) );
  NOR2_X1 u5_mult_82_U2116 ( .A1(u5_mult_82_n410), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__16_) );
  NOR2_X1 u5_mult_82_U2115 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__17_) );
  NOR2_X1 u5_mult_82_U2114 ( .A1(u5_mult_82_n406), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__18_) );
  NOR2_X1 u5_mult_82_U2113 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__19_) );
  NOR2_X1 u5_mult_82_U2112 ( .A1(u5_mult_82_n445), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__1_) );
  NOR2_X1 u5_mult_82_U2111 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__20_) );
  NOR2_X1 u5_mult_82_U2110 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__21_) );
  NOR2_X1 u5_mult_82_U2109 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__22_) );
  NOR2_X1 u5_mult_82_U2108 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__23_) );
  NOR2_X1 u5_mult_82_U2107 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__24_) );
  NOR2_X1 u5_mult_82_U2106 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__25_) );
  NOR2_X1 u5_mult_82_U2105 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__26_) );
  NOR2_X1 u5_mult_82_U2104 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__27_) );
  NOR2_X1 u5_mult_82_U2103 ( .A1(u5_mult_82_n387), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__28_) );
  NOR2_X1 u5_mult_82_U2102 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__29_) );
  NOR2_X1 u5_mult_82_U2101 ( .A1(u5_mult_82_n442), .A2(u5_mult_82_n328), .ZN(
        u5_mult_82_ab_2__2_) );
  NOR2_X1 u5_mult_82_U2100 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n328), .ZN(
        u5_mult_82_ab_2__30_) );
  NOR2_X1 u5_mult_82_U2099 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n328), .ZN(
        u5_mult_82_ab_2__31_) );
  NOR2_X1 u5_mult_82_U2098 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n328), .ZN(
        u5_mult_82_ab_2__32_) );
  NOR2_X1 u5_mult_82_U2097 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n328), .ZN(
        u5_mult_82_ab_2__33_) );
  NOR2_X1 u5_mult_82_U2096 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n328), .ZN(
        u5_mult_82_ab_2__34_) );
  NOR2_X1 u5_mult_82_U2095 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n328), .ZN(
        u5_mult_82_ab_2__35_) );
  NOR2_X1 u5_mult_82_U2094 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n328), .ZN(
        u5_mult_82_ab_2__36_) );
  NOR2_X1 u5_mult_82_U2093 ( .A1(u5_mult_82_n370), .A2(u5_mult_82_n328), .ZN(
        u5_mult_82_ab_2__37_) );
  NOR2_X1 u5_mult_82_U2092 ( .A1(u5_mult_82_n367), .A2(u5_mult_82_n328), .ZN(
        u5_mult_82_ab_2__38_) );
  NOR2_X1 u5_mult_82_U2091 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n328), .ZN(
        u5_mult_82_ab_2__39_) );
  NOR2_X1 u5_mult_82_U2090 ( .A1(u5_mult_82_n441), .A2(u5_mult_82_n329), .ZN(
        u5_mult_82_ab_2__3_) );
  NOR2_X1 u5_mult_82_U2089 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n329), .ZN(
        u5_mult_82_ab_2__40_) );
  NOR2_X1 u5_mult_82_U2088 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n329), .ZN(
        u5_mult_82_ab_2__41_) );
  NOR2_X1 u5_mult_82_U2087 ( .A1(u5_mult_82_n358), .A2(u5_mult_82_n329), .ZN(
        u5_mult_82_ab_2__42_) );
  NOR2_X1 u5_mult_82_U2086 ( .A1(u5_mult_82_n356), .A2(u5_mult_82_n329), .ZN(
        u5_mult_82_ab_2__43_) );
  NOR2_X1 u5_mult_82_U2085 ( .A1(u5_mult_82_n353), .A2(u5_mult_82_n329), .ZN(
        u5_mult_82_ab_2__44_) );
  NOR2_X1 u5_mult_82_U2084 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n329), .ZN(
        u5_mult_82_ab_2__45_) );
  NOR2_X1 u5_mult_82_U2083 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n329), .ZN(
        u5_mult_82_ab_2__46_) );
  NOR2_X1 u5_mult_82_U2082 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n329), .ZN(
        u5_mult_82_ab_2__47_) );
  NOR2_X1 u5_mult_82_U2081 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n329), .ZN(
        u5_mult_82_ab_2__48_) );
  NOR2_X1 u5_mult_82_U2080 ( .A1(u5_mult_82_n343), .A2(u5_mult_82_n329), .ZN(
        u5_mult_82_ab_2__49_) );
  NOR2_X1 u5_mult_82_U2079 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__4_) );
  NOR2_X1 u5_mult_82_U2078 ( .A1(u5_mult_82_n342), .A2(u5_mult_82_n329), .ZN(
        u5_mult_82_ab_2__50_) );
  NOR2_X1 u5_mult_82_U2077 ( .A1(u5_mult_82_n338), .A2(u5_mult_82_n328), .ZN(
        u5_mult_82_ab_2__51_) );
  NOR2_X1 u5_mult_82_U2076 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n328), .ZN(
        u5_mult_82_ab_2__52_) );
  NOR2_X1 u5_mult_82_U2075 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__5_) );
  NOR2_X1 u5_mult_82_U2074 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__6_) );
  NOR2_X1 u5_mult_82_U2073 ( .A1(u5_mult_82_n432), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__7_) );
  NOR2_X1 u5_mult_82_U2072 ( .A1(u5_mult_82_n430), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__8_) );
  NOR2_X1 u5_mult_82_U2071 ( .A1(u5_mult_82_n428), .A2(u5_mult_82_n327), .ZN(
        u5_mult_82_ab_2__9_) );
  NOR2_X1 u5_mult_82_U2070 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n270), .ZN(
        u5_mult_82_ab_30__0_) );
  NOR2_X1 u5_mult_82_U2069 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n271), .ZN(
        u5_mult_82_ab_30__10_) );
  NOR2_X1 u5_mult_82_U2068 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n270), .ZN(
        u5_mult_82_ab_30__11_) );
  NOR2_X1 u5_mult_82_U2067 ( .A1(u5_mult_82_n422), .A2(u5_mult_82_n271), .ZN(
        u5_mult_82_ab_30__12_) );
  NOR2_X1 u5_mult_82_U2066 ( .A1(u5_mult_82_n419), .A2(u5_mult_82_n270), .ZN(
        u5_mult_82_ab_30__13_) );
  NOR2_X1 u5_mult_82_U2065 ( .A1(u5_mult_82_n416), .A2(u5_mult_82_n270), .ZN(
        u5_mult_82_ab_30__14_) );
  NOR2_X1 u5_mult_82_U2064 ( .A1(u5_mult_82_n413), .A2(u5_mult_82_n270), .ZN(
        u5_mult_82_ab_30__15_) );
  NOR2_X1 u5_mult_82_U2063 ( .A1(u5_mult_82_n410), .A2(u5_mult_82_n270), .ZN(
        u5_mult_82_ab_30__16_) );
  NOR2_X1 u5_mult_82_U2062 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n270), .ZN(
        u5_mult_82_ab_30__17_) );
  NOR2_X1 u5_mult_82_U2061 ( .A1(u5_mult_82_n406), .A2(u5_mult_82_n271), .ZN(
        u5_mult_82_ab_30__18_) );
  NOR2_X1 u5_mult_82_U2060 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n271), .ZN(
        u5_mult_82_ab_30__19_) );
  NOR2_X1 u5_mult_82_U2059 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n460), .ZN(
        u5_mult_82_ab_30__1_) );
  NOR2_X1 u5_mult_82_U2058 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n460), .ZN(
        u5_mult_82_ab_30__20_) );
  NOR2_X1 u5_mult_82_U2057 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n460), .ZN(
        u5_mult_82_ab_30__21_) );
  NOR2_X1 u5_mult_82_U2056 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n460), .ZN(
        u5_mult_82_ab_30__22_) );
  NOR2_X1 u5_mult_82_U2055 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n460), .ZN(
        u5_mult_82_ab_30__23_) );
  NOR2_X1 u5_mult_82_U2054 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n460), .ZN(
        u5_mult_82_ab_30__24_) );
  NOR2_X1 u5_mult_82_U2053 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n460), .ZN(
        u5_mult_82_ab_30__25_) );
  NOR2_X1 u5_mult_82_U2052 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n271), .ZN(
        u5_mult_82_ab_30__26_) );
  NOR2_X1 u5_mult_82_U2051 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n460), .ZN(
        u5_mult_82_ab_30__27_) );
  NOR2_X1 u5_mult_82_U2050 ( .A1(u5_mult_82_n387), .A2(u5_mult_82_n460), .ZN(
        u5_mult_82_ab_30__28_) );
  NOR2_X1 u5_mult_82_U2049 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n460), .ZN(
        u5_mult_82_ab_30__29_) );
  NOR2_X1 u5_mult_82_U2048 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n270), .ZN(
        u5_mult_82_ab_30__2_) );
  NOR2_X1 u5_mult_82_U2047 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n270), .ZN(
        u5_mult_82_ab_30__30_) );
  NOR2_X1 u5_mult_82_U2046 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n270), .ZN(
        u5_mult_82_ab_30__31_) );
  NOR2_X1 u5_mult_82_U2045 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n270), .ZN(
        u5_mult_82_ab_30__32_) );
  NOR2_X1 u5_mult_82_U2044 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n270), .ZN(
        u5_mult_82_ab_30__33_) );
  NOR2_X1 u5_mult_82_U2043 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n270), .ZN(
        u5_mult_82_ab_30__34_) );
  NOR2_X1 u5_mult_82_U2042 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n270), .ZN(
        u5_mult_82_ab_30__35_) );
  NOR2_X1 u5_mult_82_U2041 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n270), .ZN(
        u5_mult_82_ab_30__36_) );
  NOR2_X1 u5_mult_82_U2040 ( .A1(u5_mult_82_n370), .A2(u5_mult_82_n270), .ZN(
        u5_mult_82_ab_30__37_) );
  NOR2_X1 u5_mult_82_U2039 ( .A1(u5_mult_82_n367), .A2(u5_mult_82_n270), .ZN(
        u5_mult_82_ab_30__38_) );
  NOR2_X1 u5_mult_82_U2038 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n270), .ZN(
        u5_mult_82_ab_30__39_) );
  NOR2_X1 u5_mult_82_U2037 ( .A1(u5_mult_82_n441), .A2(u5_mult_82_n271), .ZN(
        u5_mult_82_ab_30__3_) );
  NOR2_X1 u5_mult_82_U2036 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n271), .ZN(
        u5_mult_82_ab_30__40_) );
  NOR2_X1 u5_mult_82_U2035 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n271), .ZN(
        u5_mult_82_ab_30__41_) );
  NOR2_X1 u5_mult_82_U2034 ( .A1(u5_mult_82_n358), .A2(u5_mult_82_n271), .ZN(
        u5_mult_82_ab_30__42_) );
  NOR2_X1 u5_mult_82_U2033 ( .A1(u5_mult_82_n356), .A2(u5_mult_82_n271), .ZN(
        u5_mult_82_ab_30__43_) );
  NOR2_X1 u5_mult_82_U2032 ( .A1(u5_mult_82_n353), .A2(u5_mult_82_n271), .ZN(
        u5_mult_82_ab_30__44_) );
  NOR2_X1 u5_mult_82_U2031 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n271), .ZN(
        u5_mult_82_ab_30__45_) );
  NOR2_X1 u5_mult_82_U2030 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n271), .ZN(
        u5_mult_82_ab_30__46_) );
  NOR2_X1 u5_mult_82_U2029 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n271), .ZN(
        u5_mult_82_ab_30__47_) );
  NOR2_X1 u5_mult_82_U2028 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n271), .ZN(
        u5_mult_82_ab_30__48_) );
  NOR2_X1 u5_mult_82_U2027 ( .A1(u5_mult_82_n343), .A2(u5_mult_82_n271), .ZN(
        u5_mult_82_ab_30__49_) );
  NOR2_X1 u5_mult_82_U2026 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n270), .ZN(
        u5_mult_82_ab_30__4_) );
  NOR2_X1 u5_mult_82_U2025 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n270), .ZN(
        u5_mult_82_ab_30__50_) );
  NOR2_X1 u5_mult_82_U2024 ( .A1(u5_mult_82_n338), .A2(u5_mult_82_n270), .ZN(
        u5_mult_82_ab_30__51_) );
  NOR2_X1 u5_mult_82_U2023 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n270), .ZN(
        u5_mult_82_ab_30__52_) );
  NOR2_X1 u5_mult_82_U2022 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n270), .ZN(
        u5_mult_82_ab_30__5_) );
  NOR2_X1 u5_mult_82_U2021 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n270), .ZN(
        u5_mult_82_ab_30__6_) );
  NOR2_X1 u5_mult_82_U2020 ( .A1(u5_mult_82_n432), .A2(u5_mult_82_n270), .ZN(
        u5_mult_82_ab_30__7_) );
  NOR2_X1 u5_mult_82_U2019 ( .A1(u5_mult_82_n430), .A2(u5_mult_82_n270), .ZN(
        u5_mult_82_ab_30__8_) );
  NOR2_X1 u5_mult_82_U2018 ( .A1(u5_mult_82_n428), .A2(u5_mult_82_n271), .ZN(
        u5_mult_82_ab_30__9_) );
  NOR2_X1 u5_mult_82_U2017 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n269), .ZN(
        u5_mult_82_ab_31__0_) );
  NOR2_X1 u5_mult_82_U2016 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n269), .ZN(
        u5_mult_82_ab_31__10_) );
  NOR2_X1 u5_mult_82_U2015 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n269), .ZN(
        u5_mult_82_ab_31__11_) );
  NOR2_X1 u5_mult_82_U2014 ( .A1(u5_mult_82_n422), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__12_) );
  NOR2_X1 u5_mult_82_U2013 ( .A1(u5_mult_82_n419), .A2(u5_mult_82_n269), .ZN(
        u5_mult_82_ab_31__13_) );
  NOR2_X1 u5_mult_82_U2012 ( .A1(u5_mult_82_n416), .A2(u5_mult_82_n269), .ZN(
        u5_mult_82_ab_31__14_) );
  NOR2_X1 u5_mult_82_U2011 ( .A1(u5_mult_82_n413), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__15_) );
  NOR2_X1 u5_mult_82_U2010 ( .A1(u5_mult_82_n410), .A2(u5_mult_82_n269), .ZN(
        u5_mult_82_ab_31__16_) );
  NOR2_X1 u5_mult_82_U2009 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n269), .ZN(
        u5_mult_82_ab_31__17_) );
  NOR2_X1 u5_mult_82_U2008 ( .A1(u5_mult_82_n406), .A2(u5_mult_82_n269), .ZN(
        u5_mult_82_ab_31__18_) );
  NOR2_X1 u5_mult_82_U2007 ( .A1(u5_mult_82_n404), .A2(u5_mult_82_n269), .ZN(
        u5_mult_82_ab_31__19_) );
  NOR2_X1 u5_mult_82_U2006 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__1_) );
  NOR2_X1 u5_mult_82_U2005 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n459), .ZN(
        u5_mult_82_ab_31__20_) );
  NOR2_X1 u5_mult_82_U2004 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n459), .ZN(
        u5_mult_82_ab_31__21_) );
  NOR2_X1 u5_mult_82_U2003 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n459), .ZN(
        u5_mult_82_ab_31__22_) );
  NOR2_X1 u5_mult_82_U2002 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n459), .ZN(
        u5_mult_82_ab_31__23_) );
  NOR2_X1 u5_mult_82_U2001 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n459), .ZN(
        u5_mult_82_ab_31__24_) );
  NOR2_X1 u5_mult_82_U2000 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n459), .ZN(
        u5_mult_82_ab_31__25_) );
  NOR2_X1 u5_mult_82_U1999 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__26_) );
  NOR2_X1 u5_mult_82_U1998 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__27_) );
  NOR2_X1 u5_mult_82_U1997 ( .A1(u5_mult_82_n387), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__28_) );
  NOR2_X1 u5_mult_82_U1996 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__29_) );
  NOR2_X1 u5_mult_82_U1995 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__2_) );
  NOR2_X1 u5_mult_82_U1994 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__30_) );
  NOR2_X1 u5_mult_82_U1993 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__31_) );
  NOR2_X1 u5_mult_82_U1992 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__32_) );
  NOR2_X1 u5_mult_82_U1991 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__33_) );
  NOR2_X1 u5_mult_82_U1990 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__34_) );
  NOR2_X1 u5_mult_82_U1989 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__35_) );
  NOR2_X1 u5_mult_82_U1988 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__36_) );
  NOR2_X1 u5_mult_82_U1987 ( .A1(u5_mult_82_n370), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__37_) );
  NOR2_X1 u5_mult_82_U1986 ( .A1(u5_mult_82_n368), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__38_) );
  NOR2_X1 u5_mult_82_U1985 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__39_) );
  NOR2_X1 u5_mult_82_U1984 ( .A1(u5_mult_82_n441), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__3_) );
  NOR2_X1 u5_mult_82_U1983 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__40_) );
  NOR2_X1 u5_mult_82_U1982 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__41_) );
  NOR2_X1 u5_mult_82_U1981 ( .A1(u5_mult_82_n358), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__42_) );
  NOR2_X1 u5_mult_82_U1980 ( .A1(u5_mult_82_n356), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__43_) );
  NOR2_X1 u5_mult_82_U1979 ( .A1(u5_mult_82_n353), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__44_) );
  NOR2_X1 u5_mult_82_U1978 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__45_) );
  NOR2_X1 u5_mult_82_U1977 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__46_) );
  NOR2_X1 u5_mult_82_U1976 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__47_) );
  NOR2_X1 u5_mult_82_U1975 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__48_) );
  NOR2_X1 u5_mult_82_U1974 ( .A1(u5_mult_82_n343), .A2(u5_mult_82_n268), .ZN(
        u5_mult_82_ab_31__49_) );
  NOR2_X1 u5_mult_82_U1973 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n269), .ZN(
        u5_mult_82_ab_31__4_) );
  NOR2_X1 u5_mult_82_U1972 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n269), .ZN(
        u5_mult_82_ab_31__50_) );
  NOR2_X1 u5_mult_82_U1971 ( .A1(u5_mult_82_n338), .A2(u5_mult_82_n269), .ZN(
        u5_mult_82_ab_31__51_) );
  NOR2_X1 u5_mult_82_U1970 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n269), .ZN(
        u5_mult_82_ab_31__52_) );
  NOR2_X1 u5_mult_82_U1969 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n269), .ZN(
        u5_mult_82_ab_31__5_) );
  NOR2_X1 u5_mult_82_U1968 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n269), .ZN(
        u5_mult_82_ab_31__6_) );
  NOR2_X1 u5_mult_82_U1967 ( .A1(u5_mult_82_n432), .A2(u5_mult_82_n269), .ZN(
        u5_mult_82_ab_31__7_) );
  NOR2_X1 u5_mult_82_U1966 ( .A1(u5_mult_82_n430), .A2(u5_mult_82_n269), .ZN(
        u5_mult_82_ab_31__8_) );
  NOR2_X1 u5_mult_82_U1965 ( .A1(u5_mult_82_n428), .A2(u5_mult_82_n269), .ZN(
        u5_mult_82_ab_31__9_) );
  NOR2_X1 u5_mult_82_U1964 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n267), .ZN(
        u5_mult_82_ab_32__0_) );
  NOR2_X1 u5_mult_82_U1963 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n267), .ZN(
        u5_mult_82_ab_32__10_) );
  NOR2_X1 u5_mult_82_U1962 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n267), .ZN(
        u5_mult_82_ab_32__11_) );
  NOR2_X1 u5_mult_82_U1961 ( .A1(u5_mult_82_n422), .A2(u5_mult_82_n266), .ZN(
        u5_mult_82_ab_32__12_) );
  NOR2_X1 u5_mult_82_U1960 ( .A1(u5_mult_82_n419), .A2(u5_mult_82_n267), .ZN(
        u5_mult_82_ab_32__13_) );
  NOR2_X1 u5_mult_82_U1959 ( .A1(u5_mult_82_n416), .A2(u5_mult_82_n267), .ZN(
        u5_mult_82_ab_32__14_) );
  NOR2_X1 u5_mult_82_U1958 ( .A1(u5_mult_82_n413), .A2(u5_mult_82_n266), .ZN(
        u5_mult_82_ab_32__15_) );
  NOR2_X1 u5_mult_82_U1957 ( .A1(u5_mult_82_n410), .A2(u5_mult_82_n267), .ZN(
        u5_mult_82_ab_32__16_) );
  NOR2_X1 u5_mult_82_U1956 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n267), .ZN(
        u5_mult_82_ab_32__17_) );
  NOR2_X1 u5_mult_82_U1955 ( .A1(u5_mult_82_n406), .A2(u5_mult_82_n267), .ZN(
        u5_mult_82_ab_32__18_) );
  NOR2_X1 u5_mult_82_U1954 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n267), .ZN(
        u5_mult_82_ab_32__19_) );
  NOR2_X1 u5_mult_82_U1953 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n458), .ZN(
        u5_mult_82_ab_32__1_) );
  NOR2_X1 u5_mult_82_U1952 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n458), .ZN(
        u5_mult_82_ab_32__20_) );
  NOR2_X1 u5_mult_82_U1951 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n458), .ZN(
        u5_mult_82_ab_32__21_) );
  NOR2_X1 u5_mult_82_U1950 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n458), .ZN(
        u5_mult_82_ab_32__22_) );
  NOR2_X1 u5_mult_82_U1949 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n458), .ZN(
        u5_mult_82_ab_32__23_) );
  NOR2_X1 u5_mult_82_U1948 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n266), .ZN(
        u5_mult_82_ab_32__24_) );
  NOR2_X1 u5_mult_82_U1947 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n458), .ZN(
        u5_mult_82_ab_32__25_) );
  NOR2_X1 u5_mult_82_U1946 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n458), .ZN(
        u5_mult_82_ab_32__26_) );
  NOR2_X1 u5_mult_82_U1945 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n458), .ZN(
        u5_mult_82_ab_32__27_) );
  NOR2_X1 u5_mult_82_U1944 ( .A1(u5_mult_82_n387), .A2(u5_mult_82_n458), .ZN(
        u5_mult_82_ab_32__28_) );
  NOR2_X1 u5_mult_82_U1943 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n458), .ZN(
        u5_mult_82_ab_32__29_) );
  NOR2_X1 u5_mult_82_U1942 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n266), .ZN(
        u5_mult_82_ab_32__2_) );
  NOR2_X1 u5_mult_82_U1941 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n266), .ZN(
        u5_mult_82_ab_32__30_) );
  NOR2_X1 u5_mult_82_U1940 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n266), .ZN(
        u5_mult_82_ab_32__31_) );
  NOR2_X1 u5_mult_82_U1939 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n266), .ZN(
        u5_mult_82_ab_32__32_) );
  NOR2_X1 u5_mult_82_U1938 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n266), .ZN(
        u5_mult_82_ab_32__33_) );
  NOR2_X1 u5_mult_82_U1937 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n266), .ZN(
        u5_mult_82_ab_32__34_) );
  NOR2_X1 u5_mult_82_U1936 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n266), .ZN(
        u5_mult_82_ab_32__35_) );
  NOR2_X1 u5_mult_82_U1935 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n266), .ZN(
        u5_mult_82_ab_32__36_) );
  NOR2_X1 u5_mult_82_U1934 ( .A1(u5_mult_82_n370), .A2(u5_mult_82_n266), .ZN(
        u5_mult_82_ab_32__37_) );
  NOR2_X1 u5_mult_82_U1933 ( .A1(u5_mult_82_n367), .A2(u5_mult_82_n266), .ZN(
        u5_mult_82_ab_32__38_) );
  NOR2_X1 u5_mult_82_U1932 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n266), .ZN(
        u5_mult_82_ab_32__39_) );
  NOR2_X1 u5_mult_82_U1931 ( .A1(u5_mult_82_n440), .A2(u5_mult_82_n266), .ZN(
        u5_mult_82_ab_32__3_) );
  NOR2_X1 u5_mult_82_U1930 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n266), .ZN(
        u5_mult_82_ab_32__40_) );
  NOR2_X1 u5_mult_82_U1929 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n266), .ZN(
        u5_mult_82_ab_32__41_) );
  NOR2_X1 u5_mult_82_U1928 ( .A1(u5_mult_82_n358), .A2(u5_mult_82_n266), .ZN(
        u5_mult_82_ab_32__42_) );
  NOR2_X1 u5_mult_82_U1927 ( .A1(u5_mult_82_n356), .A2(u5_mult_82_n266), .ZN(
        u5_mult_82_ab_32__43_) );
  NOR2_X1 u5_mult_82_U1926 ( .A1(u5_mult_82_n353), .A2(u5_mult_82_n266), .ZN(
        u5_mult_82_ab_32__44_) );
  NOR2_X1 u5_mult_82_U1925 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n266), .ZN(
        u5_mult_82_ab_32__45_) );
  NOR2_X1 u5_mult_82_U1924 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n266), .ZN(
        u5_mult_82_ab_32__46_) );
  NOR2_X1 u5_mult_82_U1923 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n266), .ZN(
        u5_mult_82_ab_32__47_) );
  NOR2_X1 u5_mult_82_U1922 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n266), .ZN(
        u5_mult_82_ab_32__48_) );
  NOR2_X1 u5_mult_82_U1921 ( .A1(u5_mult_82_n343), .A2(u5_mult_82_n266), .ZN(
        u5_mult_82_ab_32__49_) );
  NOR2_X1 u5_mult_82_U1920 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n267), .ZN(
        u5_mult_82_ab_32__4_) );
  NOR2_X1 u5_mult_82_U1919 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n267), .ZN(
        u5_mult_82_ab_32__50_) );
  NOR2_X1 u5_mult_82_U1918 ( .A1(u5_mult_82_n338), .A2(u5_mult_82_n267), .ZN(
        u5_mult_82_ab_32__51_) );
  NOR2_X1 u5_mult_82_U1917 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n267), .ZN(
        u5_mult_82_ab_32__52_) );
  NOR2_X1 u5_mult_82_U1916 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n267), .ZN(
        u5_mult_82_ab_32__5_) );
  NOR2_X1 u5_mult_82_U1915 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n267), .ZN(
        u5_mult_82_ab_32__6_) );
  NOR2_X1 u5_mult_82_U1914 ( .A1(u5_mult_82_n432), .A2(u5_mult_82_n267), .ZN(
        u5_mult_82_ab_32__7_) );
  NOR2_X1 u5_mult_82_U1913 ( .A1(u5_mult_82_n430), .A2(u5_mult_82_n267), .ZN(
        u5_mult_82_ab_32__8_) );
  NOR2_X1 u5_mult_82_U1912 ( .A1(u5_mult_82_n428), .A2(u5_mult_82_n267), .ZN(
        u5_mult_82_ab_32__9_) );
  NOR2_X1 u5_mult_82_U1911 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n264), .ZN(
        u5_mult_82_ab_33__0_) );
  NOR2_X1 u5_mult_82_U1910 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n265), .ZN(
        u5_mult_82_ab_33__10_) );
  NOR2_X1 u5_mult_82_U1909 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n264), .ZN(
        u5_mult_82_ab_33__11_) );
  NOR2_X1 u5_mult_82_U1908 ( .A1(u5_mult_82_n422), .A2(u5_mult_82_n265), .ZN(
        u5_mult_82_ab_33__12_) );
  NOR2_X1 u5_mult_82_U1907 ( .A1(u5_mult_82_n419), .A2(u5_mult_82_n264), .ZN(
        u5_mult_82_ab_33__13_) );
  NOR2_X1 u5_mult_82_U1906 ( .A1(u5_mult_82_n416), .A2(u5_mult_82_n264), .ZN(
        u5_mult_82_ab_33__14_) );
  NOR2_X1 u5_mult_82_U1905 ( .A1(u5_mult_82_n413), .A2(u5_mult_82_n264), .ZN(
        u5_mult_82_ab_33__15_) );
  NOR2_X1 u5_mult_82_U1904 ( .A1(u5_mult_82_n410), .A2(u5_mult_82_n264), .ZN(
        u5_mult_82_ab_33__16_) );
  NOR2_X1 u5_mult_82_U1903 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n264), .ZN(
        u5_mult_82_ab_33__17_) );
  NOR2_X1 u5_mult_82_U1902 ( .A1(u5_mult_82_n406), .A2(u5_mult_82_n265), .ZN(
        u5_mult_82_ab_33__18_) );
  NOR2_X1 u5_mult_82_U1901 ( .A1(u5_mult_82_n404), .A2(u5_mult_82_n265), .ZN(
        u5_mult_82_ab_33__19_) );
  NOR2_X1 u5_mult_82_U1900 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n457), .ZN(
        u5_mult_82_ab_33__1_) );
  NOR2_X1 u5_mult_82_U1899 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n265), .ZN(
        u5_mult_82_ab_33__20_) );
  NOR2_X1 u5_mult_82_U1898 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n457), .ZN(
        u5_mult_82_ab_33__21_) );
  NOR2_X1 u5_mult_82_U1897 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n457), .ZN(
        u5_mult_82_ab_33__22_) );
  NOR2_X1 u5_mult_82_U1896 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n457), .ZN(
        u5_mult_82_ab_33__23_) );
  NOR2_X1 u5_mult_82_U1895 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n457), .ZN(
        u5_mult_82_ab_33__24_) );
  NOR2_X1 u5_mult_82_U1894 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n457), .ZN(
        u5_mult_82_ab_33__25_) );
  NOR2_X1 u5_mult_82_U1893 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n457), .ZN(
        u5_mult_82_ab_33__26_) );
  NOR2_X1 u5_mult_82_U1892 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n457), .ZN(
        u5_mult_82_ab_33__27_) );
  NOR2_X1 u5_mult_82_U1891 ( .A1(u5_mult_82_n387), .A2(u5_mult_82_n457), .ZN(
        u5_mult_82_ab_33__28_) );
  NOR2_X1 u5_mult_82_U1890 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n457), .ZN(
        u5_mult_82_ab_33__29_) );
  NOR2_X1 u5_mult_82_U1889 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n264), .ZN(
        u5_mult_82_ab_33__2_) );
  NOR2_X1 u5_mult_82_U1888 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n264), .ZN(
        u5_mult_82_ab_33__30_) );
  NOR2_X1 u5_mult_82_U1887 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n264), .ZN(
        u5_mult_82_ab_33__31_) );
  NOR2_X1 u5_mult_82_U1886 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n264), .ZN(
        u5_mult_82_ab_33__32_) );
  NOR2_X1 u5_mult_82_U1885 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n264), .ZN(
        u5_mult_82_ab_33__33_) );
  NOR2_X1 u5_mult_82_U1884 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n264), .ZN(
        u5_mult_82_ab_33__34_) );
  NOR2_X1 u5_mult_82_U1883 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n264), .ZN(
        u5_mult_82_ab_33__35_) );
  NOR2_X1 u5_mult_82_U1882 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n264), .ZN(
        u5_mult_82_ab_33__36_) );
  NOR2_X1 u5_mult_82_U1881 ( .A1(u5_mult_82_n370), .A2(u5_mult_82_n264), .ZN(
        u5_mult_82_ab_33__37_) );
  NOR2_X1 u5_mult_82_U1880 ( .A1(u5_mult_82_n368), .A2(u5_mult_82_n264), .ZN(
        u5_mult_82_ab_33__38_) );
  NOR2_X1 u5_mult_82_U1879 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n264), .ZN(
        u5_mult_82_ab_33__39_) );
  NOR2_X1 u5_mult_82_U1878 ( .A1(u5_mult_82_n440), .A2(u5_mult_82_n265), .ZN(
        u5_mult_82_ab_33__3_) );
  NOR2_X1 u5_mult_82_U1877 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n265), .ZN(
        u5_mult_82_ab_33__40_) );
  NOR2_X1 u5_mult_82_U1876 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n265), .ZN(
        u5_mult_82_ab_33__41_) );
  NOR2_X1 u5_mult_82_U1875 ( .A1(u5_mult_82_n358), .A2(u5_mult_82_n265), .ZN(
        u5_mult_82_ab_33__42_) );
  NOR2_X1 u5_mult_82_U1874 ( .A1(u5_mult_82_n356), .A2(u5_mult_82_n265), .ZN(
        u5_mult_82_ab_33__43_) );
  NOR2_X1 u5_mult_82_U1873 ( .A1(u5_mult_82_n353), .A2(u5_mult_82_n265), .ZN(
        u5_mult_82_ab_33__44_) );
  NOR2_X1 u5_mult_82_U1872 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n265), .ZN(
        u5_mult_82_ab_33__45_) );
  NOR2_X1 u5_mult_82_U1871 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n265), .ZN(
        u5_mult_82_ab_33__46_) );
  NOR2_X1 u5_mult_82_U1870 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n265), .ZN(
        u5_mult_82_ab_33__47_) );
  NOR2_X1 u5_mult_82_U1869 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n265), .ZN(
        u5_mult_82_ab_33__48_) );
  NOR2_X1 u5_mult_82_U1868 ( .A1(u5_mult_82_n343), .A2(u5_mult_82_n265), .ZN(
        u5_mult_82_ab_33__49_) );
  NOR2_X1 u5_mult_82_U1867 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n264), .ZN(
        u5_mult_82_ab_33__4_) );
  NOR2_X1 u5_mult_82_U1866 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n264), .ZN(
        u5_mult_82_ab_33__50_) );
  NOR2_X1 u5_mult_82_U1865 ( .A1(u5_mult_82_n338), .A2(u5_mult_82_n264), .ZN(
        u5_mult_82_ab_33__51_) );
  NOR2_X1 u5_mult_82_U1864 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n264), .ZN(
        u5_mult_82_ab_33__52_) );
  NOR2_X1 u5_mult_82_U1863 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n264), .ZN(
        u5_mult_82_ab_33__5_) );
  NOR2_X1 u5_mult_82_U1862 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n264), .ZN(
        u5_mult_82_ab_33__6_) );
  NOR2_X1 u5_mult_82_U1861 ( .A1(u5_mult_82_n432), .A2(u5_mult_82_n264), .ZN(
        u5_mult_82_ab_33__7_) );
  NOR2_X1 u5_mult_82_U1860 ( .A1(u5_mult_82_n430), .A2(u5_mult_82_n264), .ZN(
        u5_mult_82_ab_33__8_) );
  NOR2_X1 u5_mult_82_U1859 ( .A1(u5_mult_82_n428), .A2(u5_mult_82_n265), .ZN(
        u5_mult_82_ab_33__9_) );
  NOR2_X1 u5_mult_82_U1858 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n456), .ZN(
        u5_mult_82_ab_34__0_) );
  NOR2_X1 u5_mult_82_U1857 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n456), .ZN(
        u5_mult_82_ab_34__10_) );
  NOR2_X1 u5_mult_82_U1856 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n456), .ZN(
        u5_mult_82_ab_34__11_) );
  NOR2_X1 u5_mult_82_U1855 ( .A1(u5_mult_82_n422), .A2(u5_mult_82_n456), .ZN(
        u5_mult_82_ab_34__12_) );
  NOR2_X1 u5_mult_82_U1854 ( .A1(u5_mult_82_n419), .A2(u5_mult_82_n456), .ZN(
        u5_mult_82_ab_34__13_) );
  NOR2_X1 u5_mult_82_U1853 ( .A1(u5_mult_82_n416), .A2(u5_mult_82_n262), .ZN(
        u5_mult_82_ab_34__14_) );
  NOR2_X1 u5_mult_82_U1852 ( .A1(u5_mult_82_n413), .A2(u5_mult_82_n262), .ZN(
        u5_mult_82_ab_34__15_) );
  NOR2_X1 u5_mult_82_U1851 ( .A1(u5_mult_82_n410), .A2(u5_mult_82_n262), .ZN(
        u5_mult_82_ab_34__16_) );
  NOR2_X1 u5_mult_82_U1850 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n456), .ZN(
        u5_mult_82_ab_34__17_) );
  NOR2_X1 u5_mult_82_U1849 ( .A1(u5_mult_82_n406), .A2(u5_mult_82_n263), .ZN(
        u5_mult_82_ab_34__18_) );
  NOR2_X1 u5_mult_82_U1848 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n263), .ZN(
        u5_mult_82_ab_34__19_) );
  NOR2_X1 u5_mult_82_U1847 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n456), .ZN(
        u5_mult_82_ab_34__1_) );
  NOR2_X1 u5_mult_82_U1846 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n456), .ZN(
        u5_mult_82_ab_34__20_) );
  NOR2_X1 u5_mult_82_U1845 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n456), .ZN(
        u5_mult_82_ab_34__21_) );
  NOR2_X1 u5_mult_82_U1844 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n263), .ZN(
        u5_mult_82_ab_34__22_) );
  NOR2_X1 u5_mult_82_U1843 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n263), .ZN(
        u5_mult_82_ab_34__23_) );
  NOR2_X1 u5_mult_82_U1842 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n456), .ZN(
        u5_mult_82_ab_34__24_) );
  NOR2_X1 u5_mult_82_U1841 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n456), .ZN(
        u5_mult_82_ab_34__25_) );
  NOR2_X1 u5_mult_82_U1840 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n456), .ZN(
        u5_mult_82_ab_34__26_) );
  NOR2_X1 u5_mult_82_U1839 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n456), .ZN(
        u5_mult_82_ab_34__27_) );
  NOR2_X1 u5_mult_82_U1838 ( .A1(u5_mult_82_n387), .A2(u5_mult_82_n456), .ZN(
        u5_mult_82_ab_34__28_) );
  NOR2_X1 u5_mult_82_U1837 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n456), .ZN(
        u5_mult_82_ab_34__29_) );
  NOR2_X1 u5_mult_82_U1836 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n262), .ZN(
        u5_mult_82_ab_34__2_) );
  NOR2_X1 u5_mult_82_U1835 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n262), .ZN(
        u5_mult_82_ab_34__30_) );
  NOR2_X1 u5_mult_82_U1834 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n262), .ZN(
        u5_mult_82_ab_34__31_) );
  NOR2_X1 u5_mult_82_U1833 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n262), .ZN(
        u5_mult_82_ab_34__32_) );
  NOR2_X1 u5_mult_82_U1832 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n262), .ZN(
        u5_mult_82_ab_34__33_) );
  NOR2_X1 u5_mult_82_U1831 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n262), .ZN(
        u5_mult_82_ab_34__34_) );
  NOR2_X1 u5_mult_82_U1830 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n262), .ZN(
        u5_mult_82_ab_34__35_) );
  NOR2_X1 u5_mult_82_U1829 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n262), .ZN(
        u5_mult_82_ab_34__36_) );
  NOR2_X1 u5_mult_82_U1828 ( .A1(u5_mult_82_n370), .A2(u5_mult_82_n262), .ZN(
        u5_mult_82_ab_34__37_) );
  NOR2_X1 u5_mult_82_U1827 ( .A1(u5_mult_82_n367), .A2(u5_mult_82_n262), .ZN(
        u5_mult_82_ab_34__38_) );
  NOR2_X1 u5_mult_82_U1826 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n262), .ZN(
        u5_mult_82_ab_34__39_) );
  NOR2_X1 u5_mult_82_U1825 ( .A1(u5_mult_82_n440), .A2(u5_mult_82_n263), .ZN(
        u5_mult_82_ab_34__3_) );
  NOR2_X1 u5_mult_82_U1824 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n263), .ZN(
        u5_mult_82_ab_34__40_) );
  NOR2_X1 u5_mult_82_U1823 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n263), .ZN(
        u5_mult_82_ab_34__41_) );
  NOR2_X1 u5_mult_82_U1822 ( .A1(u5_mult_82_n358), .A2(u5_mult_82_n263), .ZN(
        u5_mult_82_ab_34__42_) );
  NOR2_X1 u5_mult_82_U1821 ( .A1(u5_mult_82_n356), .A2(u5_mult_82_n263), .ZN(
        u5_mult_82_ab_34__43_) );
  NOR2_X1 u5_mult_82_U1820 ( .A1(u5_mult_82_n353), .A2(u5_mult_82_n263), .ZN(
        u5_mult_82_ab_34__44_) );
  NOR2_X1 u5_mult_82_U1819 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n263), .ZN(
        u5_mult_82_ab_34__45_) );
  NOR2_X1 u5_mult_82_U1818 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n263), .ZN(
        u5_mult_82_ab_34__46_) );
  NOR2_X1 u5_mult_82_U1817 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n263), .ZN(
        u5_mult_82_ab_34__47_) );
  NOR2_X1 u5_mult_82_U1816 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n263), .ZN(
        u5_mult_82_ab_34__48_) );
  NOR2_X1 u5_mult_82_U1815 ( .A1(u5_mult_82_n343), .A2(u5_mult_82_n263), .ZN(
        u5_mult_82_ab_34__49_) );
  NOR2_X1 u5_mult_82_U1814 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n262), .ZN(
        u5_mult_82_ab_34__4_) );
  NOR2_X1 u5_mult_82_U1813 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n262), .ZN(
        u5_mult_82_ab_34__50_) );
  NOR2_X1 u5_mult_82_U1812 ( .A1(u5_mult_82_n338), .A2(u5_mult_82_n262), .ZN(
        u5_mult_82_ab_34__51_) );
  NOR2_X1 u5_mult_82_U1811 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n262), .ZN(
        u5_mult_82_ab_34__52_) );
  NOR2_X1 u5_mult_82_U1810 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n262), .ZN(
        u5_mult_82_ab_34__5_) );
  NOR2_X1 u5_mult_82_U1809 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n262), .ZN(
        u5_mult_82_ab_34__6_) );
  NOR2_X1 u5_mult_82_U1808 ( .A1(u5_mult_82_n432), .A2(u5_mult_82_n262), .ZN(
        u5_mult_82_ab_34__7_) );
  NOR2_X1 u5_mult_82_U1807 ( .A1(u5_mult_82_n430), .A2(u5_mult_82_n262), .ZN(
        u5_mult_82_ab_34__8_) );
  NOR2_X1 u5_mult_82_U1806 ( .A1(u5_mult_82_n428), .A2(u5_mult_82_n263), .ZN(
        u5_mult_82_ab_34__9_) );
  NOR2_X1 u5_mult_82_U1805 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n261), .ZN(
        u5_mult_82_ab_35__0_) );
  NOR2_X1 u5_mult_82_U1804 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n261), .ZN(
        u5_mult_82_ab_35__10_) );
  NOR2_X1 u5_mult_82_U1803 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n261), .ZN(
        u5_mult_82_ab_35__11_) );
  NOR2_X1 u5_mult_82_U1802 ( .A1(u5_mult_82_n422), .A2(u5_mult_82_n261), .ZN(
        u5_mult_82_ab_35__12_) );
  NOR2_X1 u5_mult_82_U1801 ( .A1(u5_mult_82_n419), .A2(u5_mult_82_n261), .ZN(
        u5_mult_82_ab_35__13_) );
  NOR2_X1 u5_mult_82_U1800 ( .A1(u5_mult_82_n416), .A2(u5_mult_82_n259), .ZN(
        u5_mult_82_ab_35__14_) );
  NOR2_X1 u5_mult_82_U1799 ( .A1(u5_mult_82_n413), .A2(u5_mult_82_n259), .ZN(
        u5_mult_82_ab_35__15_) );
  NOR2_X1 u5_mult_82_U1798 ( .A1(u5_mult_82_n410), .A2(u5_mult_82_n260), .ZN(
        u5_mult_82_ab_35__16_) );
  NOR2_X1 u5_mult_82_U1797 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n261), .ZN(
        u5_mult_82_ab_35__17_) );
  NOR2_X1 u5_mult_82_U1796 ( .A1(u5_mult_82_n406), .A2(u5_mult_82_n261), .ZN(
        u5_mult_82_ab_35__18_) );
  NOR2_X1 u5_mult_82_U1795 ( .A1(u5_mult_82_n404), .A2(u5_mult_82_n261), .ZN(
        u5_mult_82_ab_35__19_) );
  NOR2_X1 u5_mult_82_U1794 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n261), .ZN(
        u5_mult_82_ab_35__1_) );
  NOR2_X1 u5_mult_82_U1793 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n261), .ZN(
        u5_mult_82_ab_35__20_) );
  NOR2_X1 u5_mult_82_U1792 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n260), .ZN(
        u5_mult_82_ab_35__21_) );
  NOR2_X1 u5_mult_82_U1791 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n260), .ZN(
        u5_mult_82_ab_35__22_) );
  NOR2_X1 u5_mult_82_U1790 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n260), .ZN(
        u5_mult_82_ab_35__23_) );
  NOR2_X1 u5_mult_82_U1789 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n261), .ZN(
        u5_mult_82_ab_35__24_) );
  NOR2_X1 u5_mult_82_U1788 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n261), .ZN(
        u5_mult_82_ab_35__25_) );
  NOR2_X1 u5_mult_82_U1787 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n261), .ZN(
        u5_mult_82_ab_35__26_) );
  NOR2_X1 u5_mult_82_U1786 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n261), .ZN(
        u5_mult_82_ab_35__27_) );
  NOR2_X1 u5_mult_82_U1785 ( .A1(u5_mult_82_n387), .A2(u5_mult_82_n261), .ZN(
        u5_mult_82_ab_35__28_) );
  NOR2_X1 u5_mult_82_U1784 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n261), .ZN(
        u5_mult_82_ab_35__29_) );
  NOR2_X1 u5_mult_82_U1783 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n259), .ZN(
        u5_mult_82_ab_35__2_) );
  NOR2_X1 u5_mult_82_U1782 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n259), .ZN(
        u5_mult_82_ab_35__30_) );
  NOR2_X1 u5_mult_82_U1781 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n259), .ZN(
        u5_mult_82_ab_35__31_) );
  NOR2_X1 u5_mult_82_U1780 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n259), .ZN(
        u5_mult_82_ab_35__32_) );
  NOR2_X1 u5_mult_82_U1779 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n259), .ZN(
        u5_mult_82_ab_35__33_) );
  NOR2_X1 u5_mult_82_U1778 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n259), .ZN(
        u5_mult_82_ab_35__34_) );
  NOR2_X1 u5_mult_82_U1777 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n259), .ZN(
        u5_mult_82_ab_35__35_) );
  NOR2_X1 u5_mult_82_U1776 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n259), .ZN(
        u5_mult_82_ab_35__36_) );
  NOR2_X1 u5_mult_82_U1775 ( .A1(u5_mult_82_n370), .A2(u5_mult_82_n259), .ZN(
        u5_mult_82_ab_35__37_) );
  NOR2_X1 u5_mult_82_U1774 ( .A1(u5_mult_82_n368), .A2(u5_mult_82_n259), .ZN(
        u5_mult_82_ab_35__38_) );
  NOR2_X1 u5_mult_82_U1773 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n259), .ZN(
        u5_mult_82_ab_35__39_) );
  NOR2_X1 u5_mult_82_U1772 ( .A1(u5_mult_82_n440), .A2(u5_mult_82_n260), .ZN(
        u5_mult_82_ab_35__3_) );
  NOR2_X1 u5_mult_82_U1771 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n260), .ZN(
        u5_mult_82_ab_35__40_) );
  NOR2_X1 u5_mult_82_U1770 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n260), .ZN(
        u5_mult_82_ab_35__41_) );
  NOR2_X1 u5_mult_82_U1769 ( .A1(u5_mult_82_n358), .A2(u5_mult_82_n260), .ZN(
        u5_mult_82_ab_35__42_) );
  NOR2_X1 u5_mult_82_U1768 ( .A1(u5_mult_82_n356), .A2(u5_mult_82_n260), .ZN(
        u5_mult_82_ab_35__43_) );
  NOR2_X1 u5_mult_82_U1767 ( .A1(u5_mult_82_n353), .A2(u5_mult_82_n260), .ZN(
        u5_mult_82_ab_35__44_) );
  NOR2_X1 u5_mult_82_U1766 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n260), .ZN(
        u5_mult_82_ab_35__45_) );
  NOR2_X1 u5_mult_82_U1765 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n260), .ZN(
        u5_mult_82_ab_35__46_) );
  NOR2_X1 u5_mult_82_U1764 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n260), .ZN(
        u5_mult_82_ab_35__47_) );
  NOR2_X1 u5_mult_82_U1763 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n260), .ZN(
        u5_mult_82_ab_35__48_) );
  NOR2_X1 u5_mult_82_U1762 ( .A1(u5_mult_82_n343), .A2(u5_mult_82_n260), .ZN(
        u5_mult_82_ab_35__49_) );
  NOR2_X1 u5_mult_82_U1761 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n259), .ZN(
        u5_mult_82_ab_35__4_) );
  NOR2_X1 u5_mult_82_U1760 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n259), .ZN(
        u5_mult_82_ab_35__50_) );
  NOR2_X1 u5_mult_82_U1759 ( .A1(u5_mult_82_n338), .A2(u5_mult_82_n259), .ZN(
        u5_mult_82_ab_35__51_) );
  NOR2_X1 u5_mult_82_U1758 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n259), .ZN(
        u5_mult_82_ab_35__52_) );
  NOR2_X1 u5_mult_82_U1757 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n259), .ZN(
        u5_mult_82_ab_35__5_) );
  NOR2_X1 u5_mult_82_U1756 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n259), .ZN(
        u5_mult_82_ab_35__6_) );
  NOR2_X1 u5_mult_82_U1755 ( .A1(u5_mult_82_n432), .A2(u5_mult_82_n259), .ZN(
        u5_mult_82_ab_35__7_) );
  NOR2_X1 u5_mult_82_U1754 ( .A1(u5_mult_82_n430), .A2(u5_mult_82_n259), .ZN(
        u5_mult_82_ab_35__8_) );
  NOR2_X1 u5_mult_82_U1753 ( .A1(u5_mult_82_n428), .A2(u5_mult_82_n260), .ZN(
        u5_mult_82_ab_35__9_) );
  NOR2_X1 u5_mult_82_U1752 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n258), .ZN(
        u5_mult_82_ab_36__0_) );
  NOR2_X1 u5_mult_82_U1751 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n256), .ZN(
        u5_mult_82_ab_36__10_) );
  NOR2_X1 u5_mult_82_U1750 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n256), .ZN(
        u5_mult_82_ab_36__11_) );
  NOR2_X1 u5_mult_82_U1749 ( .A1(u5_mult_82_n422), .A2(u5_mult_82_n256), .ZN(
        u5_mult_82_ab_36__12_) );
  NOR2_X1 u5_mult_82_U1748 ( .A1(u5_mult_82_n419), .A2(u5_mult_82_n257), .ZN(
        u5_mult_82_ab_36__13_) );
  NOR2_X1 u5_mult_82_U1747 ( .A1(u5_mult_82_n416), .A2(u5_mult_82_n257), .ZN(
        u5_mult_82_ab_36__14_) );
  NOR2_X1 u5_mult_82_U1746 ( .A1(u5_mult_82_n413), .A2(u5_mult_82_n257), .ZN(
        u5_mult_82_ab_36__15_) );
  NOR2_X1 u5_mult_82_U1745 ( .A1(u5_mult_82_n410), .A2(u5_mult_82_n258), .ZN(
        u5_mult_82_ab_36__16_) );
  NOR2_X1 u5_mult_82_U1744 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n258), .ZN(
        u5_mult_82_ab_36__17_) );
  NOR2_X1 u5_mult_82_U1743 ( .A1(u5_mult_82_n406), .A2(u5_mult_82_n258), .ZN(
        u5_mult_82_ab_36__18_) );
  NOR2_X1 u5_mult_82_U1742 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n258), .ZN(
        u5_mult_82_ab_36__19_) );
  NOR2_X1 u5_mult_82_U1741 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n258), .ZN(
        u5_mult_82_ab_36__1_) );
  NOR2_X1 u5_mult_82_U1740 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n257), .ZN(
        u5_mult_82_ab_36__20_) );
  NOR2_X1 u5_mult_82_U1739 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n258), .ZN(
        u5_mult_82_ab_36__21_) );
  NOR2_X1 u5_mult_82_U1738 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n258), .ZN(
        u5_mult_82_ab_36__22_) );
  NOR2_X1 u5_mult_82_U1737 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n258), .ZN(
        u5_mult_82_ab_36__23_) );
  NOR2_X1 u5_mult_82_U1736 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n258), .ZN(
        u5_mult_82_ab_36__24_) );
  NOR2_X1 u5_mult_82_U1735 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n258), .ZN(
        u5_mult_82_ab_36__25_) );
  NOR2_X1 u5_mult_82_U1734 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n258), .ZN(
        u5_mult_82_ab_36__26_) );
  NOR2_X1 u5_mult_82_U1733 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n258), .ZN(
        u5_mult_82_ab_36__27_) );
  NOR2_X1 u5_mult_82_U1732 ( .A1(u5_mult_82_n387), .A2(u5_mult_82_n258), .ZN(
        u5_mult_82_ab_36__28_) );
  NOR2_X1 u5_mult_82_U1731 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n258), .ZN(
        u5_mult_82_ab_36__29_) );
  NOR2_X1 u5_mult_82_U1730 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n256), .ZN(
        u5_mult_82_ab_36__2_) );
  NOR2_X1 u5_mult_82_U1729 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n256), .ZN(
        u5_mult_82_ab_36__30_) );
  NOR2_X1 u5_mult_82_U1728 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n256), .ZN(
        u5_mult_82_ab_36__31_) );
  NOR2_X1 u5_mult_82_U1727 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n256), .ZN(
        u5_mult_82_ab_36__32_) );
  NOR2_X1 u5_mult_82_U1726 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n256), .ZN(
        u5_mult_82_ab_36__33_) );
  NOR2_X1 u5_mult_82_U1725 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n256), .ZN(
        u5_mult_82_ab_36__34_) );
  NOR2_X1 u5_mult_82_U1724 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n256), .ZN(
        u5_mult_82_ab_36__35_) );
  NOR2_X1 u5_mult_82_U1723 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n256), .ZN(
        u5_mult_82_ab_36__36_) );
  NOR2_X1 u5_mult_82_U1722 ( .A1(u5_mult_82_n370), .A2(u5_mult_82_n256), .ZN(
        u5_mult_82_ab_36__37_) );
  NOR2_X1 u5_mult_82_U1721 ( .A1(u5_mult_82_n367), .A2(u5_mult_82_n256), .ZN(
        u5_mult_82_ab_36__38_) );
  NOR2_X1 u5_mult_82_U1720 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n256), .ZN(
        u5_mult_82_ab_36__39_) );
  NOR2_X1 u5_mult_82_U1719 ( .A1(u5_mult_82_n441), .A2(u5_mult_82_n257), .ZN(
        u5_mult_82_ab_36__3_) );
  NOR2_X1 u5_mult_82_U1718 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n257), .ZN(
        u5_mult_82_ab_36__40_) );
  NOR2_X1 u5_mult_82_U1717 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n257), .ZN(
        u5_mult_82_ab_36__41_) );
  NOR2_X1 u5_mult_82_U1716 ( .A1(u5_mult_82_n358), .A2(u5_mult_82_n257), .ZN(
        u5_mult_82_ab_36__42_) );
  NOR2_X1 u5_mult_82_U1715 ( .A1(u5_mult_82_n356), .A2(u5_mult_82_n257), .ZN(
        u5_mult_82_ab_36__43_) );
  NOR2_X1 u5_mult_82_U1714 ( .A1(u5_mult_82_n353), .A2(u5_mult_82_n257), .ZN(
        u5_mult_82_ab_36__44_) );
  NOR2_X1 u5_mult_82_U1713 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n257), .ZN(
        u5_mult_82_ab_36__45_) );
  NOR2_X1 u5_mult_82_U1712 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n257), .ZN(
        u5_mult_82_ab_36__46_) );
  NOR2_X1 u5_mult_82_U1711 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n257), .ZN(
        u5_mult_82_ab_36__47_) );
  NOR2_X1 u5_mult_82_U1710 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n257), .ZN(
        u5_mult_82_ab_36__48_) );
  NOR2_X1 u5_mult_82_U1709 ( .A1(u5_mult_82_n343), .A2(u5_mult_82_n257), .ZN(
        u5_mult_82_ab_36__49_) );
  NOR2_X1 u5_mult_82_U1708 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n256), .ZN(
        u5_mult_82_ab_36__4_) );
  NOR2_X1 u5_mult_82_U1707 ( .A1(u5_mult_82_n342), .A2(u5_mult_82_n256), .ZN(
        u5_mult_82_ab_36__50_) );
  NOR2_X1 u5_mult_82_U1706 ( .A1(u5_mult_82_n338), .A2(u5_mult_82_n256), .ZN(
        u5_mult_82_ab_36__51_) );
  NOR2_X1 u5_mult_82_U1705 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n256), .ZN(
        u5_mult_82_ab_36__52_) );
  NOR2_X1 u5_mult_82_U1704 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n256), .ZN(
        u5_mult_82_ab_36__5_) );
  NOR2_X1 u5_mult_82_U1703 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n256), .ZN(
        u5_mult_82_ab_36__6_) );
  NOR2_X1 u5_mult_82_U1702 ( .A1(u5_mult_82_n432), .A2(u5_mult_82_n256), .ZN(
        u5_mult_82_ab_36__7_) );
  NOR2_X1 u5_mult_82_U1701 ( .A1(u5_mult_82_n430), .A2(u5_mult_82_n256), .ZN(
        u5_mult_82_ab_36__8_) );
  NOR2_X1 u5_mult_82_U1700 ( .A1(u5_mult_82_n428), .A2(u5_mult_82_n257), .ZN(
        u5_mult_82_ab_36__9_) );
  NOR2_X1 u5_mult_82_U1699 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n255), .ZN(
        u5_mult_82_ab_37__0_) );
  NOR2_X1 u5_mult_82_U1698 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n254), .ZN(
        u5_mult_82_ab_37__10_) );
  NOR2_X1 u5_mult_82_U1697 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n254), .ZN(
        u5_mult_82_ab_37__11_) );
  NOR2_X1 u5_mult_82_U1696 ( .A1(u5_mult_82_n422), .A2(u5_mult_82_n254), .ZN(
        u5_mult_82_ab_37__12_) );
  NOR2_X1 u5_mult_82_U1695 ( .A1(u5_mult_82_n419), .A2(u5_mult_82_n255), .ZN(
        u5_mult_82_ab_37__13_) );
  NOR2_X1 u5_mult_82_U1694 ( .A1(u5_mult_82_n416), .A2(u5_mult_82_n253), .ZN(
        u5_mult_82_ab_37__14_) );
  NOR2_X1 u5_mult_82_U1693 ( .A1(u5_mult_82_n413), .A2(u5_mult_82_n255), .ZN(
        u5_mult_82_ab_37__15_) );
  NOR2_X1 u5_mult_82_U1692 ( .A1(u5_mult_82_n410), .A2(u5_mult_82_n253), .ZN(
        u5_mult_82_ab_37__16_) );
  NOR2_X1 u5_mult_82_U1691 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n255), .ZN(
        u5_mult_82_ab_37__17_) );
  NOR2_X1 u5_mult_82_U1690 ( .A1(u5_mult_82_n406), .A2(u5_mult_82_n253), .ZN(
        u5_mult_82_ab_37__18_) );
  NOR2_X1 u5_mult_82_U1689 ( .A1(u5_mult_82_n404), .A2(u5_mult_82_n253), .ZN(
        u5_mult_82_ab_37__19_) );
  NOR2_X1 u5_mult_82_U1688 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n253), .ZN(
        u5_mult_82_ab_37__1_) );
  NOR2_X1 u5_mult_82_U1687 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n253), .ZN(
        u5_mult_82_ab_37__20_) );
  NOR2_X1 u5_mult_82_U1686 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n253), .ZN(
        u5_mult_82_ab_37__21_) );
  NOR2_X1 u5_mult_82_U1685 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n253), .ZN(
        u5_mult_82_ab_37__22_) );
  NOR2_X1 u5_mult_82_U1684 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n253), .ZN(
        u5_mult_82_ab_37__23_) );
  NOR2_X1 u5_mult_82_U1683 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n253), .ZN(
        u5_mult_82_ab_37__24_) );
  NOR2_X1 u5_mult_82_U1682 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n253), .ZN(
        u5_mult_82_ab_37__25_) );
  NOR2_X1 u5_mult_82_U1681 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n253), .ZN(
        u5_mult_82_ab_37__26_) );
  NOR2_X1 u5_mult_82_U1680 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n253), .ZN(
        u5_mult_82_ab_37__27_) );
  NOR2_X1 u5_mult_82_U1679 ( .A1(u5_mult_82_n387), .A2(u5_mult_82_n253), .ZN(
        u5_mult_82_ab_37__28_) );
  NOR2_X1 u5_mult_82_U1678 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n253), .ZN(
        u5_mult_82_ab_37__29_) );
  NOR2_X1 u5_mult_82_U1677 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n254), .ZN(
        u5_mult_82_ab_37__2_) );
  NOR2_X1 u5_mult_82_U1676 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n254), .ZN(
        u5_mult_82_ab_37__30_) );
  NOR2_X1 u5_mult_82_U1675 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n254), .ZN(
        u5_mult_82_ab_37__31_) );
  NOR2_X1 u5_mult_82_U1674 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n254), .ZN(
        u5_mult_82_ab_37__32_) );
  NOR2_X1 u5_mult_82_U1673 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n254), .ZN(
        u5_mult_82_ab_37__33_) );
  NOR2_X1 u5_mult_82_U1672 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n254), .ZN(
        u5_mult_82_ab_37__34_) );
  NOR2_X1 u5_mult_82_U1671 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n254), .ZN(
        u5_mult_82_ab_37__35_) );
  NOR2_X1 u5_mult_82_U1670 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n254), .ZN(
        u5_mult_82_ab_37__36_) );
  NOR2_X1 u5_mult_82_U1669 ( .A1(u5_mult_82_n370), .A2(u5_mult_82_n254), .ZN(
        u5_mult_82_ab_37__37_) );
  NOR2_X1 u5_mult_82_U1668 ( .A1(u5_mult_82_n368), .A2(u5_mult_82_n254), .ZN(
        u5_mult_82_ab_37__38_) );
  NOR2_X1 u5_mult_82_U1667 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n254), .ZN(
        u5_mult_82_ab_37__39_) );
  NOR2_X1 u5_mult_82_U1666 ( .A1(u5_mult_82_n478), .A2(u5_mult_82_n255), .ZN(
        u5_mult_82_ab_37__3_) );
  NOR2_X1 u5_mult_82_U1665 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n255), .ZN(
        u5_mult_82_ab_37__40_) );
  NOR2_X1 u5_mult_82_U1664 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n255), .ZN(
        u5_mult_82_ab_37__41_) );
  NOR2_X1 u5_mult_82_U1663 ( .A1(u5_mult_82_n358), .A2(u5_mult_82_n255), .ZN(
        u5_mult_82_ab_37__42_) );
  NOR2_X1 u5_mult_82_U1662 ( .A1(u5_mult_82_n356), .A2(u5_mult_82_n255), .ZN(
        u5_mult_82_ab_37__43_) );
  NOR2_X1 u5_mult_82_U1661 ( .A1(u5_mult_82_n353), .A2(u5_mult_82_n255), .ZN(
        u5_mult_82_ab_37__44_) );
  NOR2_X1 u5_mult_82_U1660 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n255), .ZN(
        u5_mult_82_ab_37__45_) );
  NOR2_X1 u5_mult_82_U1659 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n255), .ZN(
        u5_mult_82_ab_37__46_) );
  NOR2_X1 u5_mult_82_U1658 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n255), .ZN(
        u5_mult_82_ab_37__47_) );
  NOR2_X1 u5_mult_82_U1657 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n255), .ZN(
        u5_mult_82_ab_37__48_) );
  NOR2_X1 u5_mult_82_U1656 ( .A1(u5_mult_82_n343), .A2(u5_mult_82_n255), .ZN(
        u5_mult_82_ab_37__49_) );
  NOR2_X1 u5_mult_82_U1655 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n254), .ZN(
        u5_mult_82_ab_37__4_) );
  NOR2_X1 u5_mult_82_U1654 ( .A1(u5_mult_82_n342), .A2(u5_mult_82_n254), .ZN(
        u5_mult_82_ab_37__50_) );
  NOR2_X1 u5_mult_82_U1653 ( .A1(u5_mult_82_n338), .A2(u5_mult_82_n254), .ZN(
        u5_mult_82_ab_37__51_) );
  NOR2_X1 u5_mult_82_U1652 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n254), .ZN(
        u5_mult_82_ab_37__52_) );
  NOR2_X1 u5_mult_82_U1651 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n254), .ZN(
        u5_mult_82_ab_37__5_) );
  NOR2_X1 u5_mult_82_U1650 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n254), .ZN(
        u5_mult_82_ab_37__6_) );
  NOR2_X1 u5_mult_82_U1649 ( .A1(u5_mult_82_n432), .A2(u5_mult_82_n254), .ZN(
        u5_mult_82_ab_37__7_) );
  NOR2_X1 u5_mult_82_U1648 ( .A1(u5_mult_82_n430), .A2(u5_mult_82_n255), .ZN(
        u5_mult_82_ab_37__8_) );
  NOR2_X1 u5_mult_82_U1647 ( .A1(u5_mult_82_n428), .A2(u5_mult_82_n253), .ZN(
        u5_mult_82_ab_37__9_) );
  NOR2_X1 u5_mult_82_U1646 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n250), .ZN(
        u5_mult_82_ab_38__0_) );
  NOR2_X1 u5_mult_82_U1645 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n250), .ZN(
        u5_mult_82_ab_38__10_) );
  NOR2_X1 u5_mult_82_U1644 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n251), .ZN(
        u5_mult_82_ab_38__11_) );
  NOR2_X1 u5_mult_82_U1643 ( .A1(u5_mult_82_n422), .A2(u5_mult_82_n249), .ZN(
        u5_mult_82_ab_38__12_) );
  NOR2_X1 u5_mult_82_U1642 ( .A1(u5_mult_82_n419), .A2(u5_mult_82_n252), .ZN(
        u5_mult_82_ab_38__13_) );
  NOR2_X1 u5_mult_82_U1641 ( .A1(u5_mult_82_n416), .A2(u5_mult_82_n252), .ZN(
        u5_mult_82_ab_38__14_) );
  NOR2_X1 u5_mult_82_U1640 ( .A1(u5_mult_82_n413), .A2(u5_mult_82_n252), .ZN(
        u5_mult_82_ab_38__15_) );
  NOR2_X1 u5_mult_82_U1639 ( .A1(u5_mult_82_n410), .A2(u5_mult_82_n252), .ZN(
        u5_mult_82_ab_38__16_) );
  NOR2_X1 u5_mult_82_U1638 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n252), .ZN(
        u5_mult_82_ab_38__17_) );
  NOR2_X1 u5_mult_82_U1637 ( .A1(u5_mult_82_n406), .A2(u5_mult_82_n249), .ZN(
        u5_mult_82_ab_38__18_) );
  NOR2_X1 u5_mult_82_U1636 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n250), .ZN(
        u5_mult_82_ab_38__19_) );
  NOR2_X1 u5_mult_82_U1635 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n249), .ZN(
        u5_mult_82_ab_38__1_) );
  NOR2_X1 u5_mult_82_U1634 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n249), .ZN(
        u5_mult_82_ab_38__20_) );
  NOR2_X1 u5_mult_82_U1633 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n249), .ZN(
        u5_mult_82_ab_38__21_) );
  NOR2_X1 u5_mult_82_U1632 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n249), .ZN(
        u5_mult_82_ab_38__22_) );
  NOR2_X1 u5_mult_82_U1631 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n249), .ZN(
        u5_mult_82_ab_38__23_) );
  NOR2_X1 u5_mult_82_U1630 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n249), .ZN(
        u5_mult_82_ab_38__24_) );
  NOR2_X1 u5_mult_82_U1629 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n249), .ZN(
        u5_mult_82_ab_38__25_) );
  NOR2_X1 u5_mult_82_U1628 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n249), .ZN(
        u5_mult_82_ab_38__26_) );
  NOR2_X1 u5_mult_82_U1627 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n249), .ZN(
        u5_mult_82_ab_38__27_) );
  NOR2_X1 u5_mult_82_U1626 ( .A1(u5_mult_82_n387), .A2(u5_mult_82_n249), .ZN(
        u5_mult_82_ab_38__28_) );
  NOR2_X1 u5_mult_82_U1625 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n249), .ZN(
        u5_mult_82_ab_38__29_) );
  NOR2_X1 u5_mult_82_U1624 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n250), .ZN(
        u5_mult_82_ab_38__2_) );
  NOR2_X1 u5_mult_82_U1623 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n250), .ZN(
        u5_mult_82_ab_38__30_) );
  NOR2_X1 u5_mult_82_U1622 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n250), .ZN(
        u5_mult_82_ab_38__31_) );
  NOR2_X1 u5_mult_82_U1621 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n250), .ZN(
        u5_mult_82_ab_38__32_) );
  NOR2_X1 u5_mult_82_U1620 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n250), .ZN(
        u5_mult_82_ab_38__33_) );
  NOR2_X1 u5_mult_82_U1619 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n250), .ZN(
        u5_mult_82_ab_38__34_) );
  NOR2_X1 u5_mult_82_U1618 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n250), .ZN(
        u5_mult_82_ab_38__35_) );
  NOR2_X1 u5_mult_82_U1617 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n250), .ZN(
        u5_mult_82_ab_38__36_) );
  NOR2_X1 u5_mult_82_U1616 ( .A1(u5_mult_82_n370), .A2(u5_mult_82_n250), .ZN(
        u5_mult_82_ab_38__37_) );
  NOR2_X1 u5_mult_82_U1615 ( .A1(u5_mult_82_n369), .A2(u5_mult_82_n250), .ZN(
        u5_mult_82_ab_38__38_) );
  NOR2_X1 u5_mult_82_U1614 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n250), .ZN(
        u5_mult_82_ab_38__39_) );
  NOR2_X1 u5_mult_82_U1613 ( .A1(u5_mult_82_n478), .A2(u5_mult_82_n251), .ZN(
        u5_mult_82_ab_38__3_) );
  NOR2_X1 u5_mult_82_U1612 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n251), .ZN(
        u5_mult_82_ab_38__40_) );
  NOR2_X1 u5_mult_82_U1611 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n251), .ZN(
        u5_mult_82_ab_38__41_) );
  NOR2_X1 u5_mult_82_U1610 ( .A1(u5_mult_82_n358), .A2(u5_mult_82_n251), .ZN(
        u5_mult_82_ab_38__42_) );
  NOR2_X1 u5_mult_82_U1609 ( .A1(u5_mult_82_n356), .A2(u5_mult_82_n251), .ZN(
        u5_mult_82_ab_38__43_) );
  NOR2_X1 u5_mult_82_U1608 ( .A1(u5_mult_82_n353), .A2(u5_mult_82_n251), .ZN(
        u5_mult_82_ab_38__44_) );
  NOR2_X1 u5_mult_82_U1607 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n251), .ZN(
        u5_mult_82_ab_38__45_) );
  NOR2_X1 u5_mult_82_U1606 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n251), .ZN(
        u5_mult_82_ab_38__46_) );
  NOR2_X1 u5_mult_82_U1605 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n251), .ZN(
        u5_mult_82_ab_38__47_) );
  NOR2_X1 u5_mult_82_U1604 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n251), .ZN(
        u5_mult_82_ab_38__48_) );
  NOR2_X1 u5_mult_82_U1603 ( .A1(u5_mult_82_n343), .A2(u5_mult_82_n251), .ZN(
        u5_mult_82_ab_38__49_) );
  NOR2_X1 u5_mult_82_U1602 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n250), .ZN(
        u5_mult_82_ab_38__4_) );
  NOR2_X1 u5_mult_82_U1601 ( .A1(u5_mult_82_n342), .A2(u5_mult_82_n250), .ZN(
        u5_mult_82_ab_38__50_) );
  NOR2_X1 u5_mult_82_U1600 ( .A1(u5_mult_82_n338), .A2(u5_mult_82_n250), .ZN(
        u5_mult_82_ab_38__51_) );
  NOR2_X1 u5_mult_82_U1599 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n250), .ZN(
        u5_mult_82_ab_38__52_) );
  NOR2_X1 u5_mult_82_U1598 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n250), .ZN(
        u5_mult_82_ab_38__5_) );
  NOR2_X1 u5_mult_82_U1597 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n250), .ZN(
        u5_mult_82_ab_38__6_) );
  NOR2_X1 u5_mult_82_U1596 ( .A1(u5_mult_82_n432), .A2(u5_mult_82_n250), .ZN(
        u5_mult_82_ab_38__7_) );
  NOR2_X1 u5_mult_82_U1595 ( .A1(u5_mult_82_n430), .A2(u5_mult_82_n249), .ZN(
        u5_mult_82_ab_38__8_) );
  NOR2_X1 u5_mult_82_U1594 ( .A1(u5_mult_82_n428), .A2(u5_mult_82_n251), .ZN(
        u5_mult_82_ab_38__9_) );
  NOR2_X1 u5_mult_82_U1593 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__0_) );
  NOR2_X1 u5_mult_82_U1592 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n248), .ZN(
        u5_mult_82_ab_39__10_) );
  NOR2_X1 u5_mult_82_U1591 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n455), .ZN(
        u5_mult_82_ab_39__11_) );
  NOR2_X1 u5_mult_82_U1590 ( .A1(u5_mult_82_n422), .A2(u5_mult_82_n455), .ZN(
        u5_mult_82_ab_39__12_) );
  NOR2_X1 u5_mult_82_U1589 ( .A1(u5_mult_82_n419), .A2(u5_mult_82_n455), .ZN(
        u5_mult_82_ab_39__13_) );
  NOR2_X1 u5_mult_82_U1588 ( .A1(u5_mult_82_n416), .A2(u5_mult_82_n455), .ZN(
        u5_mult_82_ab_39__14_) );
  NOR2_X1 u5_mult_82_U1587 ( .A1(u5_mult_82_n413), .A2(u5_mult_82_n455), .ZN(
        u5_mult_82_ab_39__15_) );
  NOR2_X1 u5_mult_82_U1586 ( .A1(u5_mult_82_n410), .A2(u5_mult_82_n455), .ZN(
        u5_mult_82_ab_39__16_) );
  NOR2_X1 u5_mult_82_U1585 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n248), .ZN(
        u5_mult_82_ab_39__17_) );
  NOR2_X1 u5_mult_82_U1584 ( .A1(u5_mult_82_n406), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__18_) );
  NOR2_X1 u5_mult_82_U1583 ( .A1(u5_mult_82_n404), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__19_) );
  NOR2_X1 u5_mult_82_U1582 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__1_) );
  NOR2_X1 u5_mult_82_U1581 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__20_) );
  NOR2_X1 u5_mult_82_U1580 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__21_) );
  NOR2_X1 u5_mult_82_U1579 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__22_) );
  NOR2_X1 u5_mult_82_U1578 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__23_) );
  NOR2_X1 u5_mult_82_U1577 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__24_) );
  NOR2_X1 u5_mult_82_U1576 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__25_) );
  NOR2_X1 u5_mult_82_U1575 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__26_) );
  NOR2_X1 u5_mult_82_U1574 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__27_) );
  NOR2_X1 u5_mult_82_U1573 ( .A1(u5_mult_82_n387), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__28_) );
  NOR2_X1 u5_mult_82_U1572 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__29_) );
  NOR2_X1 u5_mult_82_U1571 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__2_) );
  NOR2_X1 u5_mult_82_U1570 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__30_) );
  NOR2_X1 u5_mult_82_U1569 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__31_) );
  NOR2_X1 u5_mult_82_U1568 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__32_) );
  NOR2_X1 u5_mult_82_U1567 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__33_) );
  NOR2_X1 u5_mult_82_U1566 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__34_) );
  NOR2_X1 u5_mult_82_U1565 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__35_) );
  NOR2_X1 u5_mult_82_U1564 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__36_) );
  NOR2_X1 u5_mult_82_U1563 ( .A1(u5_mult_82_n370), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__37_) );
  NOR2_X1 u5_mult_82_U1562 ( .A1(u5_mult_82_n369), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__38_) );
  NOR2_X1 u5_mult_82_U1561 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__39_) );
  NOR2_X1 u5_mult_82_U1560 ( .A1(u5_mult_82_n478), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__3_) );
  NOR2_X1 u5_mult_82_U1559 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__40_) );
  NOR2_X1 u5_mult_82_U1558 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__41_) );
  NOR2_X1 u5_mult_82_U1557 ( .A1(u5_mult_82_n358), .A2(u5_mult_82_n248), .ZN(
        u5_mult_82_ab_39__42_) );
  NOR2_X1 u5_mult_82_U1556 ( .A1(u5_mult_82_n356), .A2(u5_mult_82_n248), .ZN(
        u5_mult_82_ab_39__43_) );
  NOR2_X1 u5_mult_82_U1555 ( .A1(u5_mult_82_n353), .A2(u5_mult_82_n248), .ZN(
        u5_mult_82_ab_39__44_) );
  NOR2_X1 u5_mult_82_U1554 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__45_) );
  NOR2_X1 u5_mult_82_U1553 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n248), .ZN(
        u5_mult_82_ab_39__46_) );
  NOR2_X1 u5_mult_82_U1552 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n248), .ZN(
        u5_mult_82_ab_39__47_) );
  NOR2_X1 u5_mult_82_U1551 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n248), .ZN(
        u5_mult_82_ab_39__48_) );
  NOR2_X1 u5_mult_82_U1550 ( .A1(u5_mult_82_n343), .A2(u5_mult_82_n247), .ZN(
        u5_mult_82_ab_39__49_) );
  NOR2_X1 u5_mult_82_U1549 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n248), .ZN(
        u5_mult_82_ab_39__4_) );
  NOR2_X1 u5_mult_82_U1548 ( .A1(u5_mult_82_n342), .A2(u5_mult_82_n248), .ZN(
        u5_mult_82_ab_39__50_) );
  NOR2_X1 u5_mult_82_U1547 ( .A1(u5_mult_82_n338), .A2(u5_mult_82_n248), .ZN(
        u5_mult_82_ab_39__51_) );
  NOR2_X1 u5_mult_82_U1546 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n248), .ZN(
        u5_mult_82_ab_39__52_) );
  NOR2_X1 u5_mult_82_U1545 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n248), .ZN(
        u5_mult_82_ab_39__5_) );
  NOR2_X1 u5_mult_82_U1544 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n248), .ZN(
        u5_mult_82_ab_39__6_) );
  NOR2_X1 u5_mult_82_U1543 ( .A1(u5_mult_82_n432), .A2(u5_mult_82_n248), .ZN(
        u5_mult_82_ab_39__7_) );
  NOR2_X1 u5_mult_82_U1542 ( .A1(u5_mult_82_n430), .A2(u5_mult_82_n248), .ZN(
        u5_mult_82_ab_39__8_) );
  NOR2_X1 u5_mult_82_U1541 ( .A1(u5_mult_82_n428), .A2(u5_mult_82_n248), .ZN(
        u5_mult_82_ab_39__9_) );
  NOR2_X1 u5_mult_82_U1540 ( .A1(u5_mult_82_n480), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__0_) );
  NOR2_X1 u5_mult_82_U1539 ( .A1(u5_mult_82_n477), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__10_) );
  NOR2_X1 u5_mult_82_U1538 ( .A1(u5_mult_82_n426), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__11_) );
  NOR2_X1 u5_mult_82_U1537 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__12_) );
  NOR2_X1 u5_mult_82_U1536 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__13_) );
  NOR2_X1 u5_mult_82_U1535 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__14_) );
  NOR2_X1 u5_mult_82_U1534 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__15_) );
  NOR2_X1 u5_mult_82_U1533 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__16_) );
  NOR2_X1 u5_mult_82_U1532 ( .A1(u5_mult_82_n409), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__17_) );
  NOR2_X1 u5_mult_82_U1531 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__18_) );
  NOR2_X1 u5_mult_82_U1530 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__19_) );
  NOR2_X1 u5_mult_82_U1529 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__1_) );
  NOR2_X1 u5_mult_82_U1528 ( .A1(u5_mult_82_n475), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__20_) );
  NOR2_X1 u5_mult_82_U1527 ( .A1(u5_mult_82_n402), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__21_) );
  NOR2_X1 u5_mult_82_U1526 ( .A1(u5_mult_82_n400), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__22_) );
  NOR2_X1 u5_mult_82_U1525 ( .A1(u5_mult_82_n398), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__23_) );
  NOR2_X1 u5_mult_82_U1524 ( .A1(u5_mult_82_n396), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__24_) );
  NOR2_X1 u5_mult_82_U1523 ( .A1(u5_mult_82_n394), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__25_) );
  NOR2_X1 u5_mult_82_U1522 ( .A1(u5_mult_82_n392), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__26_) );
  NOR2_X1 u5_mult_82_U1521 ( .A1(u5_mult_82_n390), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__27_) );
  NOR2_X1 u5_mult_82_U1520 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__28_) );
  NOR2_X1 u5_mult_82_U1519 ( .A1(u5_mult_82_n386), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__29_) );
  NOR2_X1 u5_mult_82_U1518 ( .A1(u5_mult_82_n442), .A2(u5_mult_82_n326), .ZN(
        u5_mult_82_ab_3__2_) );
  NOR2_X1 u5_mult_82_U1517 ( .A1(u5_mult_82_n384), .A2(u5_mult_82_n326), .ZN(
        u5_mult_82_ab_3__30_) );
  NOR2_X1 u5_mult_82_U1516 ( .A1(u5_mult_82_n382), .A2(u5_mult_82_n326), .ZN(
        u5_mult_82_ab_3__31_) );
  NOR2_X1 u5_mult_82_U1515 ( .A1(u5_mult_82_n380), .A2(u5_mult_82_n326), .ZN(
        u5_mult_82_ab_3__32_) );
  NOR2_X1 u5_mult_82_U1514 ( .A1(u5_mult_82_n378), .A2(u5_mult_82_n326), .ZN(
        u5_mult_82_ab_3__33_) );
  NOR2_X1 u5_mult_82_U1513 ( .A1(u5_mult_82_n376), .A2(u5_mult_82_n326), .ZN(
        u5_mult_82_ab_3__34_) );
  NOR2_X1 u5_mult_82_U1512 ( .A1(u5_mult_82_n374), .A2(u5_mult_82_n326), .ZN(
        u5_mult_82_ab_3__35_) );
  NOR2_X1 u5_mult_82_U1511 ( .A1(u5_mult_82_n474), .A2(u5_mult_82_n326), .ZN(
        u5_mult_82_ab_3__36_) );
  NOR2_X1 u5_mult_82_U1510 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n326), .ZN(
        u5_mult_82_ab_3__37_) );
  NOR2_X1 u5_mult_82_U1509 ( .A1(u5_mult_82_n367), .A2(u5_mult_82_n326), .ZN(
        u5_mult_82_ab_3__38_) );
  NOR2_X1 u5_mult_82_U1508 ( .A1(u5_mult_82_n366), .A2(u5_mult_82_n326), .ZN(
        u5_mult_82_ab_3__39_) );
  NOR2_X1 u5_mult_82_U1507 ( .A1(u5_mult_82_n441), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__3_) );
  NOR2_X1 u5_mult_82_U1506 ( .A1(u5_mult_82_n364), .A2(u5_mult_82_n326), .ZN(
        u5_mult_82_ab_3__40_) );
  NOR2_X1 u5_mult_82_U1505 ( .A1(u5_mult_82_n362), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__41_) );
  NOR2_X1 u5_mult_82_U1504 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__42_) );
  NOR2_X1 u5_mult_82_U1503 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__43_) );
  NOR2_X1 u5_mult_82_U1502 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__44_) );
  NOR2_X1 u5_mult_82_U1501 ( .A1(u5_mult_82_n352), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__45_) );
  NOR2_X1 u5_mult_82_U1500 ( .A1(u5_mult_82_n350), .A2(u5_mult_82_n326), .ZN(
        u5_mult_82_ab_3__46_) );
  NOR2_X1 u5_mult_82_U1499 ( .A1(u5_mult_82_n348), .A2(u5_mult_82_n326), .ZN(
        u5_mult_82_ab_3__47_) );
  NOR2_X1 u5_mult_82_U1498 ( .A1(u5_mult_82_n346), .A2(u5_mult_82_n326), .ZN(
        u5_mult_82_ab_3__48_) );
  NOR2_X1 u5_mult_82_U1497 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n326), .ZN(
        u5_mult_82_ab_3__49_) );
  NOR2_X1 u5_mult_82_U1496 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__4_) );
  NOR2_X1 u5_mult_82_U1495 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n326), .ZN(
        u5_mult_82_ab_3__50_) );
  NOR2_X1 u5_mult_82_U1494 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n326), .ZN(
        u5_mult_82_ab_3__51_) );
  NOR2_X1 u5_mult_82_U1493 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n326), .ZN(
        u5_mult_82_ab_3__52_) );
  NOR2_X1 u5_mult_82_U1492 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__5_) );
  NOR2_X1 u5_mult_82_U1491 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__6_) );
  NOR2_X1 u5_mult_82_U1490 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__7_) );
  NOR2_X1 u5_mult_82_U1489 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__8_) );
  NOR2_X1 u5_mult_82_U1488 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n325), .ZN(
        u5_mult_82_ab_3__9_) );
  NOR2_X1 u5_mult_82_U1487 ( .A1(u5_mult_82_n480), .A2(u5_mult_82_n244), .ZN(
        u5_mult_82_ab_40__0_) );
  NOR2_X1 u5_mult_82_U1486 ( .A1(u5_mult_82_n477), .A2(u5_mult_82_n245), .ZN(
        u5_mult_82_ab_40__10_) );
  NOR2_X1 u5_mult_82_U1485 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n246), .ZN(
        u5_mult_82_ab_40__11_) );
  NOR2_X1 u5_mult_82_U1484 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n245), .ZN(
        u5_mult_82_ab_40__12_) );
  NOR2_X1 u5_mult_82_U1483 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n245), .ZN(
        u5_mult_82_ab_40__13_) );
  NOR2_X1 u5_mult_82_U1482 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n246), .ZN(
        u5_mult_82_ab_40__14_) );
  NOR2_X1 u5_mult_82_U1481 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n246), .ZN(
        u5_mult_82_ab_40__15_) );
  NOR2_X1 u5_mult_82_U1480 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n245), .ZN(
        u5_mult_82_ab_40__16_) );
  NOR2_X1 u5_mult_82_U1479 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n244), .ZN(
        u5_mult_82_ab_40__17_) );
  NOR2_X1 u5_mult_82_U1478 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n244), .ZN(
        u5_mult_82_ab_40__18_) );
  NOR2_X1 u5_mult_82_U1477 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n244), .ZN(
        u5_mult_82_ab_40__19_) );
  NOR2_X1 u5_mult_82_U1476 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n244), .ZN(
        u5_mult_82_ab_40__1_) );
  NOR2_X1 u5_mult_82_U1475 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n244), .ZN(
        u5_mult_82_ab_40__20_) );
  NOR2_X1 u5_mult_82_U1474 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n244), .ZN(
        u5_mult_82_ab_40__21_) );
  NOR2_X1 u5_mult_82_U1473 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n244), .ZN(
        u5_mult_82_ab_40__22_) );
  NOR2_X1 u5_mult_82_U1472 ( .A1(u5_mult_82_n398), .A2(u5_mult_82_n244), .ZN(
        u5_mult_82_ab_40__23_) );
  NOR2_X1 u5_mult_82_U1471 ( .A1(u5_mult_82_n396), .A2(u5_mult_82_n244), .ZN(
        u5_mult_82_ab_40__24_) );
  NOR2_X1 u5_mult_82_U1470 ( .A1(u5_mult_82_n394), .A2(u5_mult_82_n244), .ZN(
        u5_mult_82_ab_40__25_) );
  NOR2_X1 u5_mult_82_U1469 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n244), .ZN(
        u5_mult_82_ab_40__26_) );
  NOR2_X1 u5_mult_82_U1468 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n244), .ZN(
        u5_mult_82_ab_40__27_) );
  NOR2_X1 u5_mult_82_U1467 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n244), .ZN(
        u5_mult_82_ab_40__28_) );
  NOR2_X1 u5_mult_82_U1466 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n244), .ZN(
        u5_mult_82_ab_40__29_) );
  NOR2_X1 u5_mult_82_U1465 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n245), .ZN(
        u5_mult_82_ab_40__2_) );
  NOR2_X1 u5_mult_82_U1464 ( .A1(u5_mult_82_n384), .A2(u5_mult_82_n245), .ZN(
        u5_mult_82_ab_40__30_) );
  NOR2_X1 u5_mult_82_U1463 ( .A1(u5_mult_82_n382), .A2(u5_mult_82_n245), .ZN(
        u5_mult_82_ab_40__31_) );
  NOR2_X1 u5_mult_82_U1462 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n245), .ZN(
        u5_mult_82_ab_40__32_) );
  NOR2_X1 u5_mult_82_U1461 ( .A1(u5_mult_82_n378), .A2(u5_mult_82_n245), .ZN(
        u5_mult_82_ab_40__33_) );
  NOR2_X1 u5_mult_82_U1460 ( .A1(u5_mult_82_n376), .A2(u5_mult_82_n245), .ZN(
        u5_mult_82_ab_40__34_) );
  NOR2_X1 u5_mult_82_U1459 ( .A1(u5_mult_82_n374), .A2(u5_mult_82_n245), .ZN(
        u5_mult_82_ab_40__35_) );
  NOR2_X1 u5_mult_82_U1458 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n245), .ZN(
        u5_mult_82_ab_40__36_) );
  NOR2_X1 u5_mult_82_U1457 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n245), .ZN(
        u5_mult_82_ab_40__37_) );
  NOR2_X1 u5_mult_82_U1456 ( .A1(u5_mult_82_n367), .A2(u5_mult_82_n245), .ZN(
        u5_mult_82_ab_40__38_) );
  NOR2_X1 u5_mult_82_U1455 ( .A1(u5_mult_82_n366), .A2(u5_mult_82_n245), .ZN(
        u5_mult_82_ab_40__39_) );
  NOR2_X1 u5_mult_82_U1454 ( .A1(u5_mult_82_n478), .A2(u5_mult_82_n246), .ZN(
        u5_mult_82_ab_40__3_) );
  NOR2_X1 u5_mult_82_U1453 ( .A1(u5_mult_82_n364), .A2(u5_mult_82_n246), .ZN(
        u5_mult_82_ab_40__40_) );
  NOR2_X1 u5_mult_82_U1452 ( .A1(u5_mult_82_n362), .A2(u5_mult_82_n246), .ZN(
        u5_mult_82_ab_40__41_) );
  NOR2_X1 u5_mult_82_U1451 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n246), .ZN(
        u5_mult_82_ab_40__42_) );
  NOR2_X1 u5_mult_82_U1450 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n246), .ZN(
        u5_mult_82_ab_40__43_) );
  NOR2_X1 u5_mult_82_U1449 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n246), .ZN(
        u5_mult_82_ab_40__44_) );
  NOR2_X1 u5_mult_82_U1448 ( .A1(u5_mult_82_n352), .A2(u5_mult_82_n246), .ZN(
        u5_mult_82_ab_40__45_) );
  NOR2_X1 u5_mult_82_U1447 ( .A1(u5_mult_82_n350), .A2(u5_mult_82_n246), .ZN(
        u5_mult_82_ab_40__46_) );
  NOR2_X1 u5_mult_82_U1446 ( .A1(u5_mult_82_n348), .A2(u5_mult_82_n246), .ZN(
        u5_mult_82_ab_40__47_) );
  NOR2_X1 u5_mult_82_U1445 ( .A1(u5_mult_82_n346), .A2(u5_mult_82_n246), .ZN(
        u5_mult_82_ab_40__48_) );
  NOR2_X1 u5_mult_82_U1444 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n246), .ZN(
        u5_mult_82_ab_40__49_) );
  NOR2_X1 u5_mult_82_U1443 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n244), .ZN(
        u5_mult_82_ab_40__4_) );
  NOR2_X1 u5_mult_82_U1442 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n244), .ZN(
        u5_mult_82_ab_40__50_) );
  NOR2_X1 u5_mult_82_U1441 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n244), .ZN(
        u5_mult_82_ab_40__51_) );
  NOR2_X1 u5_mult_82_U1440 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n244), .ZN(
        u5_mult_82_ab_40__52_) );
  NOR2_X1 u5_mult_82_U1439 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n244), .ZN(
        u5_mult_82_ab_40__5_) );
  NOR2_X1 u5_mult_82_U1438 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n244), .ZN(
        u5_mult_82_ab_40__6_) );
  NOR2_X1 u5_mult_82_U1437 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n244), .ZN(
        u5_mult_82_ab_40__7_) );
  NOR2_X1 u5_mult_82_U1436 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n245), .ZN(
        u5_mult_82_ab_40__8_) );
  NOR2_X1 u5_mult_82_U1435 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n246), .ZN(
        u5_mult_82_ab_40__9_) );
  NOR2_X1 u5_mult_82_U1434 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n242), .ZN(
        u5_mult_82_ab_41__0_) );
  NOR2_X1 u5_mult_82_U1433 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n243), .ZN(
        u5_mult_82_ab_41__10_) );
  NOR2_X1 u5_mult_82_U1432 ( .A1(u5_mult_82_n426), .A2(u5_mult_82_n243), .ZN(
        u5_mult_82_ab_41__11_) );
  NOR2_X1 u5_mult_82_U1431 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n243), .ZN(
        u5_mult_82_ab_41__12_) );
  NOR2_X1 u5_mult_82_U1430 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n243), .ZN(
        u5_mult_82_ab_41__13_) );
  NOR2_X1 u5_mult_82_U1429 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n243), .ZN(
        u5_mult_82_ab_41__14_) );
  NOR2_X1 u5_mult_82_U1428 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n241), .ZN(
        u5_mult_82_ab_41__15_) );
  NOR2_X1 u5_mult_82_U1427 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n240), .ZN(
        u5_mult_82_ab_41__16_) );
  NOR2_X1 u5_mult_82_U1426 ( .A1(u5_mult_82_n409), .A2(u5_mult_82_n240), .ZN(
        u5_mult_82_ab_41__17_) );
  NOR2_X1 u5_mult_82_U1425 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n240), .ZN(
        u5_mult_82_ab_41__18_) );
  NOR2_X1 u5_mult_82_U1424 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n241), .ZN(
        u5_mult_82_ab_41__19_) );
  NOR2_X1 u5_mult_82_U1423 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n240), .ZN(
        u5_mult_82_ab_41__1_) );
  NOR2_X1 u5_mult_82_U1422 ( .A1(u5_mult_82_n475), .A2(u5_mult_82_n240), .ZN(
        u5_mult_82_ab_41__20_) );
  NOR2_X1 u5_mult_82_U1421 ( .A1(u5_mult_82_n402), .A2(u5_mult_82_n240), .ZN(
        u5_mult_82_ab_41__21_) );
  NOR2_X1 u5_mult_82_U1420 ( .A1(u5_mult_82_n400), .A2(u5_mult_82_n240), .ZN(
        u5_mult_82_ab_41__22_) );
  NOR2_X1 u5_mult_82_U1419 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n240), .ZN(
        u5_mult_82_ab_41__23_) );
  NOR2_X1 u5_mult_82_U1418 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n240), .ZN(
        u5_mult_82_ab_41__24_) );
  NOR2_X1 u5_mult_82_U1417 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n240), .ZN(
        u5_mult_82_ab_41__25_) );
  NOR2_X1 u5_mult_82_U1416 ( .A1(u5_mult_82_n392), .A2(u5_mult_82_n240), .ZN(
        u5_mult_82_ab_41__26_) );
  NOR2_X1 u5_mult_82_U1415 ( .A1(u5_mult_82_n390), .A2(u5_mult_82_n240), .ZN(
        u5_mult_82_ab_41__27_) );
  NOR2_X1 u5_mult_82_U1414 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n240), .ZN(
        u5_mult_82_ab_41__28_) );
  NOR2_X1 u5_mult_82_U1413 ( .A1(u5_mult_82_n386), .A2(u5_mult_82_n240), .ZN(
        u5_mult_82_ab_41__29_) );
  NOR2_X1 u5_mult_82_U1412 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n241), .ZN(
        u5_mult_82_ab_41__2_) );
  NOR2_X1 u5_mult_82_U1411 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n241), .ZN(
        u5_mult_82_ab_41__30_) );
  NOR2_X1 u5_mult_82_U1410 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n241), .ZN(
        u5_mult_82_ab_41__31_) );
  NOR2_X1 u5_mult_82_U1409 ( .A1(u5_mult_82_n380), .A2(u5_mult_82_n241), .ZN(
        u5_mult_82_ab_41__32_) );
  NOR2_X1 u5_mult_82_U1408 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n241), .ZN(
        u5_mult_82_ab_41__33_) );
  NOR2_X1 u5_mult_82_U1407 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n241), .ZN(
        u5_mult_82_ab_41__34_) );
  NOR2_X1 u5_mult_82_U1406 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n241), .ZN(
        u5_mult_82_ab_41__35_) );
  NOR2_X1 u5_mult_82_U1405 ( .A1(u5_mult_82_n474), .A2(u5_mult_82_n241), .ZN(
        u5_mult_82_ab_41__36_) );
  NOR2_X1 u5_mult_82_U1404 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n241), .ZN(
        u5_mult_82_ab_41__37_) );
  NOR2_X1 u5_mult_82_U1403 ( .A1(u5_mult_82_n367), .A2(u5_mult_82_n241), .ZN(
        u5_mult_82_ab_41__38_) );
  NOR2_X1 u5_mult_82_U1402 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n241), .ZN(
        u5_mult_82_ab_41__39_) );
  NOR2_X1 u5_mult_82_U1401 ( .A1(u5_mult_82_n478), .A2(u5_mult_82_n242), .ZN(
        u5_mult_82_ab_41__3_) );
  NOR2_X1 u5_mult_82_U1400 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n242), .ZN(
        u5_mult_82_ab_41__40_) );
  NOR2_X1 u5_mult_82_U1399 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n242), .ZN(
        u5_mult_82_ab_41__41_) );
  NOR2_X1 u5_mult_82_U1398 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n242), .ZN(
        u5_mult_82_ab_41__42_) );
  NOR2_X1 u5_mult_82_U1397 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n242), .ZN(
        u5_mult_82_ab_41__43_) );
  NOR2_X1 u5_mult_82_U1396 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n242), .ZN(
        u5_mult_82_ab_41__44_) );
  NOR2_X1 u5_mult_82_U1395 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n242), .ZN(
        u5_mult_82_ab_41__45_) );
  NOR2_X1 u5_mult_82_U1394 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n242), .ZN(
        u5_mult_82_ab_41__46_) );
  NOR2_X1 u5_mult_82_U1393 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n242), .ZN(
        u5_mult_82_ab_41__47_) );
  NOR2_X1 u5_mult_82_U1392 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n242), .ZN(
        u5_mult_82_ab_41__48_) );
  NOR2_X1 u5_mult_82_U1391 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n242), .ZN(
        u5_mult_82_ab_41__49_) );
  NOR2_X1 u5_mult_82_U1390 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n240), .ZN(
        u5_mult_82_ab_41__4_) );
  NOR2_X1 u5_mult_82_U1389 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n240), .ZN(
        u5_mult_82_ab_41__50_) );
  NOR2_X1 u5_mult_82_U1388 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n240), .ZN(
        u5_mult_82_ab_41__51_) );
  NOR2_X1 u5_mult_82_U1387 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n240), .ZN(
        u5_mult_82_ab_41__52_) );
  NOR2_X1 u5_mult_82_U1386 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n240), .ZN(
        u5_mult_82_ab_41__5_) );
  NOR2_X1 u5_mult_82_U1385 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n240), .ZN(
        u5_mult_82_ab_41__6_) );
  NOR2_X1 u5_mult_82_U1384 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n240), .ZN(
        u5_mult_82_ab_41__7_) );
  NOR2_X1 u5_mult_82_U1383 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n241), .ZN(
        u5_mult_82_ab_41__8_) );
  NOR2_X1 u5_mult_82_U1382 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n242), .ZN(
        u5_mult_82_ab_41__9_) );
  NOR2_X1 u5_mult_82_U1381 ( .A1(u5_mult_82_n480), .A2(u5_mult_82_n239), .ZN(
        u5_mult_82_ab_42__0_) );
  NOR2_X1 u5_mult_82_U1380 ( .A1(u5_mult_82_n477), .A2(u5_mult_82_n237), .ZN(
        u5_mult_82_ab_42__10_) );
  NOR2_X1 u5_mult_82_U1379 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n239), .ZN(
        u5_mult_82_ab_42__11_) );
  NOR2_X1 u5_mult_82_U1378 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n239), .ZN(
        u5_mult_82_ab_42__12_) );
  NOR2_X1 u5_mult_82_U1377 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n239), .ZN(
        u5_mult_82_ab_42__13_) );
  NOR2_X1 u5_mult_82_U1376 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n236), .ZN(
        u5_mult_82_ab_42__14_) );
  NOR2_X1 u5_mult_82_U1375 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n236), .ZN(
        u5_mult_82_ab_42__15_) );
  NOR2_X1 u5_mult_82_U1374 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n239), .ZN(
        u5_mult_82_ab_42__16_) );
  NOR2_X1 u5_mult_82_U1373 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n239), .ZN(
        u5_mult_82_ab_42__17_) );
  NOR2_X1 u5_mult_82_U1372 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n239), .ZN(
        u5_mult_82_ab_42__18_) );
  NOR2_X1 u5_mult_82_U1371 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n239), .ZN(
        u5_mult_82_ab_42__19_) );
  NOR2_X1 u5_mult_82_U1370 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n236), .ZN(
        u5_mult_82_ab_42__1_) );
  NOR2_X1 u5_mult_82_U1369 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n236), .ZN(
        u5_mult_82_ab_42__20_) );
  NOR2_X1 u5_mult_82_U1368 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n236), .ZN(
        u5_mult_82_ab_42__21_) );
  NOR2_X1 u5_mult_82_U1367 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n236), .ZN(
        u5_mult_82_ab_42__22_) );
  NOR2_X1 u5_mult_82_U1366 ( .A1(u5_mult_82_n398), .A2(u5_mult_82_n236), .ZN(
        u5_mult_82_ab_42__23_) );
  NOR2_X1 u5_mult_82_U1365 ( .A1(u5_mult_82_n396), .A2(u5_mult_82_n236), .ZN(
        u5_mult_82_ab_42__24_) );
  NOR2_X1 u5_mult_82_U1364 ( .A1(u5_mult_82_n394), .A2(u5_mult_82_n236), .ZN(
        u5_mult_82_ab_42__25_) );
  NOR2_X1 u5_mult_82_U1363 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n236), .ZN(
        u5_mult_82_ab_42__26_) );
  NOR2_X1 u5_mult_82_U1362 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n236), .ZN(
        u5_mult_82_ab_42__27_) );
  NOR2_X1 u5_mult_82_U1361 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n236), .ZN(
        u5_mult_82_ab_42__28_) );
  NOR2_X1 u5_mult_82_U1360 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n236), .ZN(
        u5_mult_82_ab_42__29_) );
  NOR2_X1 u5_mult_82_U1359 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n237), .ZN(
        u5_mult_82_ab_42__2_) );
  NOR2_X1 u5_mult_82_U1358 ( .A1(u5_mult_82_n384), .A2(u5_mult_82_n237), .ZN(
        u5_mult_82_ab_42__30_) );
  NOR2_X1 u5_mult_82_U1357 ( .A1(u5_mult_82_n382), .A2(u5_mult_82_n237), .ZN(
        u5_mult_82_ab_42__31_) );
  NOR2_X1 u5_mult_82_U1356 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n237), .ZN(
        u5_mult_82_ab_42__32_) );
  NOR2_X1 u5_mult_82_U1355 ( .A1(u5_mult_82_n378), .A2(u5_mult_82_n237), .ZN(
        u5_mult_82_ab_42__33_) );
  NOR2_X1 u5_mult_82_U1354 ( .A1(u5_mult_82_n376), .A2(u5_mult_82_n237), .ZN(
        u5_mult_82_ab_42__34_) );
  NOR2_X1 u5_mult_82_U1353 ( .A1(u5_mult_82_n374), .A2(u5_mult_82_n237), .ZN(
        u5_mult_82_ab_42__35_) );
  NOR2_X1 u5_mult_82_U1352 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n237), .ZN(
        u5_mult_82_ab_42__36_) );
  NOR2_X1 u5_mult_82_U1351 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n237), .ZN(
        u5_mult_82_ab_42__37_) );
  NOR2_X1 u5_mult_82_U1350 ( .A1(u5_mult_82_n367), .A2(u5_mult_82_n237), .ZN(
        u5_mult_82_ab_42__38_) );
  NOR2_X1 u5_mult_82_U1349 ( .A1(u5_mult_82_n366), .A2(u5_mult_82_n237), .ZN(
        u5_mult_82_ab_42__39_) );
  NOR2_X1 u5_mult_82_U1348 ( .A1(u5_mult_82_n478), .A2(u5_mult_82_n238), .ZN(
        u5_mult_82_ab_42__3_) );
  NOR2_X1 u5_mult_82_U1347 ( .A1(u5_mult_82_n364), .A2(u5_mult_82_n238), .ZN(
        u5_mult_82_ab_42__40_) );
  NOR2_X1 u5_mult_82_U1346 ( .A1(u5_mult_82_n362), .A2(u5_mult_82_n238), .ZN(
        u5_mult_82_ab_42__41_) );
  NOR2_X1 u5_mult_82_U1345 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n238), .ZN(
        u5_mult_82_ab_42__42_) );
  NOR2_X1 u5_mult_82_U1344 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n238), .ZN(
        u5_mult_82_ab_42__43_) );
  NOR2_X1 u5_mult_82_U1343 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n238), .ZN(
        u5_mult_82_ab_42__44_) );
  NOR2_X1 u5_mult_82_U1342 ( .A1(u5_mult_82_n352), .A2(u5_mult_82_n238), .ZN(
        u5_mult_82_ab_42__45_) );
  NOR2_X1 u5_mult_82_U1341 ( .A1(u5_mult_82_n350), .A2(u5_mult_82_n238), .ZN(
        u5_mult_82_ab_42__46_) );
  NOR2_X1 u5_mult_82_U1340 ( .A1(u5_mult_82_n348), .A2(u5_mult_82_n238), .ZN(
        u5_mult_82_ab_42__47_) );
  NOR2_X1 u5_mult_82_U1339 ( .A1(u5_mult_82_n346), .A2(u5_mult_82_n238), .ZN(
        u5_mult_82_ab_42__48_) );
  NOR2_X1 u5_mult_82_U1338 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n238), .ZN(
        u5_mult_82_ab_42__49_) );
  NOR2_X1 u5_mult_82_U1337 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n236), .ZN(
        u5_mult_82_ab_42__4_) );
  NOR2_X1 u5_mult_82_U1336 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n236), .ZN(
        u5_mult_82_ab_42__50_) );
  NOR2_X1 u5_mult_82_U1335 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n236), .ZN(
        u5_mult_82_ab_42__51_) );
  NOR2_X1 u5_mult_82_U1334 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n236), .ZN(
        u5_mult_82_ab_42__52_) );
  NOR2_X1 u5_mult_82_U1333 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n236), .ZN(
        u5_mult_82_ab_42__5_) );
  NOR2_X1 u5_mult_82_U1332 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n236), .ZN(
        u5_mult_82_ab_42__6_) );
  NOR2_X1 u5_mult_82_U1331 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n236), .ZN(
        u5_mult_82_ab_42__7_) );
  NOR2_X1 u5_mult_82_U1330 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n237), .ZN(
        u5_mult_82_ab_42__8_) );
  NOR2_X1 u5_mult_82_U1329 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n238), .ZN(
        u5_mult_82_ab_42__9_) );
  NOR2_X1 u5_mult_82_U1328 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n234), .ZN(
        u5_mult_82_ab_43__0_) );
  NOR2_X1 u5_mult_82_U1327 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n454), .ZN(
        u5_mult_82_ab_43__10_) );
  NOR2_X1 u5_mult_82_U1326 ( .A1(u5_mult_82_n426), .A2(u5_mult_82_n234), .ZN(
        u5_mult_82_ab_43__11_) );
  NOR2_X1 u5_mult_82_U1325 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n234), .ZN(
        u5_mult_82_ab_43__12_) );
  NOR2_X1 u5_mult_82_U1324 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n232), .ZN(
        u5_mult_82_ab_43__13_) );
  NOR2_X1 u5_mult_82_U1323 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n232), .ZN(
        u5_mult_82_ab_43__14_) );
  NOR2_X1 u5_mult_82_U1322 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n234), .ZN(
        u5_mult_82_ab_43__15_) );
  NOR2_X1 u5_mult_82_U1321 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n234), .ZN(
        u5_mult_82_ab_43__16_) );
  NOR2_X1 u5_mult_82_U1320 ( .A1(u5_mult_82_n409), .A2(u5_mult_82_n234), .ZN(
        u5_mult_82_ab_43__17_) );
  NOR2_X1 u5_mult_82_U1319 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n454), .ZN(
        u5_mult_82_ab_43__18_) );
  NOR2_X1 u5_mult_82_U1318 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n454), .ZN(
        u5_mult_82_ab_43__19_) );
  NOR2_X1 u5_mult_82_U1317 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n232), .ZN(
        u5_mult_82_ab_43__1_) );
  NOR2_X1 u5_mult_82_U1316 ( .A1(u5_mult_82_n475), .A2(u5_mult_82_n232), .ZN(
        u5_mult_82_ab_43__20_) );
  NOR2_X1 u5_mult_82_U1315 ( .A1(u5_mult_82_n402), .A2(u5_mult_82_n232), .ZN(
        u5_mult_82_ab_43__21_) );
  NOR2_X1 u5_mult_82_U1314 ( .A1(u5_mult_82_n400), .A2(u5_mult_82_n232), .ZN(
        u5_mult_82_ab_43__22_) );
  NOR2_X1 u5_mult_82_U1313 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n232), .ZN(
        u5_mult_82_ab_43__23_) );
  NOR2_X1 u5_mult_82_U1312 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n232), .ZN(
        u5_mult_82_ab_43__24_) );
  NOR2_X1 u5_mult_82_U1311 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n232), .ZN(
        u5_mult_82_ab_43__25_) );
  NOR2_X1 u5_mult_82_U1310 ( .A1(u5_mult_82_n392), .A2(u5_mult_82_n232), .ZN(
        u5_mult_82_ab_43__26_) );
  NOR2_X1 u5_mult_82_U1309 ( .A1(u5_mult_82_n390), .A2(u5_mult_82_n232), .ZN(
        u5_mult_82_ab_43__27_) );
  NOR2_X1 u5_mult_82_U1308 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n232), .ZN(
        u5_mult_82_ab_43__28_) );
  NOR2_X1 u5_mult_82_U1307 ( .A1(u5_mult_82_n386), .A2(u5_mult_82_n232), .ZN(
        u5_mult_82_ab_43__29_) );
  NOR2_X1 u5_mult_82_U1306 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n233), .ZN(
        u5_mult_82_ab_43__2_) );
  NOR2_X1 u5_mult_82_U1305 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n232), .ZN(
        u5_mult_82_ab_43__30_) );
  NOR2_X1 u5_mult_82_U1304 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n233), .ZN(
        u5_mult_82_ab_43__31_) );
  NOR2_X1 u5_mult_82_U1303 ( .A1(u5_mult_82_n380), .A2(u5_mult_82_n232), .ZN(
        u5_mult_82_ab_43__32_) );
  NOR2_X1 u5_mult_82_U1302 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n454), .ZN(
        u5_mult_82_ab_43__33_) );
  NOR2_X1 u5_mult_82_U1301 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n454), .ZN(
        u5_mult_82_ab_43__34_) );
  NOR2_X1 u5_mult_82_U1300 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n454), .ZN(
        u5_mult_82_ab_43__35_) );
  NOR2_X1 u5_mult_82_U1299 ( .A1(u5_mult_82_n474), .A2(u5_mult_82_n454), .ZN(
        u5_mult_82_ab_43__36_) );
  NOR2_X1 u5_mult_82_U1298 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n454), .ZN(
        u5_mult_82_ab_43__37_) );
  NOR2_X1 u5_mult_82_U1297 ( .A1(u5_mult_82_n367), .A2(u5_mult_82_n454), .ZN(
        u5_mult_82_ab_43__38_) );
  NOR2_X1 u5_mult_82_U1296 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n454), .ZN(
        u5_mult_82_ab_43__39_) );
  NOR2_X1 u5_mult_82_U1295 ( .A1(u5_mult_82_n441), .A2(u5_mult_82_n233), .ZN(
        u5_mult_82_ab_43__3_) );
  NOR2_X1 u5_mult_82_U1294 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n233), .ZN(
        u5_mult_82_ab_43__40_) );
  NOR2_X1 u5_mult_82_U1293 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n233), .ZN(
        u5_mult_82_ab_43__41_) );
  NOR2_X1 u5_mult_82_U1292 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n233), .ZN(
        u5_mult_82_ab_43__42_) );
  NOR2_X1 u5_mult_82_U1291 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n233), .ZN(
        u5_mult_82_ab_43__43_) );
  NOR2_X1 u5_mult_82_U1290 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n233), .ZN(
        u5_mult_82_ab_43__44_) );
  NOR2_X1 u5_mult_82_U1289 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n233), .ZN(
        u5_mult_82_ab_43__45_) );
  NOR2_X1 u5_mult_82_U1288 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n233), .ZN(
        u5_mult_82_ab_43__46_) );
  NOR2_X1 u5_mult_82_U1287 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n233), .ZN(
        u5_mult_82_ab_43__47_) );
  NOR2_X1 u5_mult_82_U1286 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n233), .ZN(
        u5_mult_82_ab_43__48_) );
  NOR2_X1 u5_mult_82_U1285 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n233), .ZN(
        u5_mult_82_ab_43__49_) );
  NOR2_X1 u5_mult_82_U1284 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n232), .ZN(
        u5_mult_82_ab_43__4_) );
  NOR2_X1 u5_mult_82_U1283 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n232), .ZN(
        u5_mult_82_ab_43__50_) );
  NOR2_X1 u5_mult_82_U1282 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n232), .ZN(
        u5_mult_82_ab_43__51_) );
  NOR2_X1 u5_mult_82_U1281 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n232), .ZN(
        u5_mult_82_ab_43__52_) );
  NOR2_X1 u5_mult_82_U1280 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n232), .ZN(
        u5_mult_82_ab_43__5_) );
  NOR2_X1 u5_mult_82_U1279 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n232), .ZN(
        u5_mult_82_ab_43__6_) );
  NOR2_X1 u5_mult_82_U1278 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n232), .ZN(
        u5_mult_82_ab_43__7_) );
  NOR2_X1 u5_mult_82_U1277 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n233), .ZN(
        u5_mult_82_ab_43__8_) );
  NOR2_X1 u5_mult_82_U1276 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n233), .ZN(
        u5_mult_82_ab_43__9_) );
  NOR2_X1 u5_mult_82_U1275 ( .A1(u5_mult_82_n480), .A2(u5_mult_82_n231), .ZN(
        u5_mult_82_ab_44__0_) );
  NOR2_X1 u5_mult_82_U1274 ( .A1(u5_mult_82_n477), .A2(u5_mult_82_n231), .ZN(
        u5_mult_82_ab_44__10_) );
  NOR2_X1 u5_mult_82_U1273 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n230), .ZN(
        u5_mult_82_ab_44__11_) );
  NOR2_X1 u5_mult_82_U1272 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n229), .ZN(
        u5_mult_82_ab_44__12_) );
  NOR2_X1 u5_mult_82_U1271 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n230), .ZN(
        u5_mult_82_ab_44__13_) );
  NOR2_X1 u5_mult_82_U1270 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n229), .ZN(
        u5_mult_82_ab_44__14_) );
  NOR2_X1 u5_mult_82_U1269 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n231), .ZN(
        u5_mult_82_ab_44__15_) );
  NOR2_X1 u5_mult_82_U1268 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n231), .ZN(
        u5_mult_82_ab_44__16_) );
  NOR2_X1 u5_mult_82_U1267 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n231), .ZN(
        u5_mult_82_ab_44__17_) );
  NOR2_X1 u5_mult_82_U1266 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n231), .ZN(
        u5_mult_82_ab_44__18_) );
  NOR2_X1 u5_mult_82_U1265 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n453), .ZN(
        u5_mult_82_ab_44__19_) );
  NOR2_X1 u5_mult_82_U1264 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n229), .ZN(
        u5_mult_82_ab_44__1_) );
  NOR2_X1 u5_mult_82_U1263 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n229), .ZN(
        u5_mult_82_ab_44__20_) );
  NOR2_X1 u5_mult_82_U1262 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n229), .ZN(
        u5_mult_82_ab_44__21_) );
  NOR2_X1 u5_mult_82_U1261 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n229), .ZN(
        u5_mult_82_ab_44__22_) );
  NOR2_X1 u5_mult_82_U1260 ( .A1(u5_mult_82_n398), .A2(u5_mult_82_n229), .ZN(
        u5_mult_82_ab_44__23_) );
  NOR2_X1 u5_mult_82_U1259 ( .A1(u5_mult_82_n396), .A2(u5_mult_82_n229), .ZN(
        u5_mult_82_ab_44__24_) );
  NOR2_X1 u5_mult_82_U1258 ( .A1(u5_mult_82_n394), .A2(u5_mult_82_n229), .ZN(
        u5_mult_82_ab_44__25_) );
  NOR2_X1 u5_mult_82_U1257 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n229), .ZN(
        u5_mult_82_ab_44__26_) );
  NOR2_X1 u5_mult_82_U1256 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n229), .ZN(
        u5_mult_82_ab_44__27_) );
  NOR2_X1 u5_mult_82_U1255 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n229), .ZN(
        u5_mult_82_ab_44__28_) );
  NOR2_X1 u5_mult_82_U1254 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n229), .ZN(
        u5_mult_82_ab_44__29_) );
  NOR2_X1 u5_mult_82_U1253 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n230), .ZN(
        u5_mult_82_ab_44__2_) );
  NOR2_X1 u5_mult_82_U1252 ( .A1(u5_mult_82_n384), .A2(u5_mult_82_n230), .ZN(
        u5_mult_82_ab_44__30_) );
  NOR2_X1 u5_mult_82_U1251 ( .A1(u5_mult_82_n382), .A2(u5_mult_82_n230), .ZN(
        u5_mult_82_ab_44__31_) );
  NOR2_X1 u5_mult_82_U1250 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n230), .ZN(
        u5_mult_82_ab_44__32_) );
  NOR2_X1 u5_mult_82_U1249 ( .A1(u5_mult_82_n378), .A2(u5_mult_82_n230), .ZN(
        u5_mult_82_ab_44__33_) );
  NOR2_X1 u5_mult_82_U1248 ( .A1(u5_mult_82_n376), .A2(u5_mult_82_n230), .ZN(
        u5_mult_82_ab_44__34_) );
  NOR2_X1 u5_mult_82_U1247 ( .A1(u5_mult_82_n374), .A2(u5_mult_82_n230), .ZN(
        u5_mult_82_ab_44__35_) );
  NOR2_X1 u5_mult_82_U1246 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n230), .ZN(
        u5_mult_82_ab_44__36_) );
  NOR2_X1 u5_mult_82_U1245 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n230), .ZN(
        u5_mult_82_ab_44__37_) );
  NOR2_X1 u5_mult_82_U1244 ( .A1(u5_mult_82_n367), .A2(u5_mult_82_n230), .ZN(
        u5_mult_82_ab_44__38_) );
  NOR2_X1 u5_mult_82_U1243 ( .A1(u5_mult_82_n366), .A2(u5_mult_82_n230), .ZN(
        u5_mult_82_ab_44__39_) );
  NOR2_X1 u5_mult_82_U1242 ( .A1(u5_mult_82_n478), .A2(u5_mult_82_n453), .ZN(
        u5_mult_82_ab_44__3_) );
  NOR2_X1 u5_mult_82_U1241 ( .A1(u5_mult_82_n364), .A2(u5_mult_82_n453), .ZN(
        u5_mult_82_ab_44__40_) );
  NOR2_X1 u5_mult_82_U1240 ( .A1(u5_mult_82_n362), .A2(u5_mult_82_n453), .ZN(
        u5_mult_82_ab_44__41_) );
  NOR2_X1 u5_mult_82_U1239 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n453), .ZN(
        u5_mult_82_ab_44__42_) );
  NOR2_X1 u5_mult_82_U1238 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n453), .ZN(
        u5_mult_82_ab_44__43_) );
  NOR2_X1 u5_mult_82_U1237 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n453), .ZN(
        u5_mult_82_ab_44__44_) );
  NOR2_X1 u5_mult_82_U1236 ( .A1(u5_mult_82_n352), .A2(u5_mult_82_n453), .ZN(
        u5_mult_82_ab_44__45_) );
  NOR2_X1 u5_mult_82_U1235 ( .A1(u5_mult_82_n350), .A2(u5_mult_82_n453), .ZN(
        u5_mult_82_ab_44__46_) );
  NOR2_X1 u5_mult_82_U1234 ( .A1(u5_mult_82_n348), .A2(u5_mult_82_n453), .ZN(
        u5_mult_82_ab_44__47_) );
  NOR2_X1 u5_mult_82_U1233 ( .A1(u5_mult_82_n346), .A2(u5_mult_82_n453), .ZN(
        u5_mult_82_ab_44__48_) );
  NOR2_X1 u5_mult_82_U1232 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n453), .ZN(
        u5_mult_82_ab_44__49_) );
  NOR2_X1 u5_mult_82_U1231 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n229), .ZN(
        u5_mult_82_ab_44__4_) );
  NOR2_X1 u5_mult_82_U1230 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n229), .ZN(
        u5_mult_82_ab_44__50_) );
  NOR2_X1 u5_mult_82_U1229 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n229), .ZN(
        u5_mult_82_ab_44__51_) );
  NOR2_X1 u5_mult_82_U1228 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n229), .ZN(
        u5_mult_82_ab_44__52_) );
  NOR2_X1 u5_mult_82_U1227 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n229), .ZN(
        u5_mult_82_ab_44__5_) );
  NOR2_X1 u5_mult_82_U1226 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n229), .ZN(
        u5_mult_82_ab_44__6_) );
  NOR2_X1 u5_mult_82_U1225 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n229), .ZN(
        u5_mult_82_ab_44__7_) );
  NOR2_X1 u5_mult_82_U1224 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n230), .ZN(
        u5_mult_82_ab_44__8_) );
  NOR2_X1 u5_mult_82_U1223 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n453), .ZN(
        u5_mult_82_ab_44__9_) );
  NOR2_X1 u5_mult_82_U1222 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n452), .ZN(
        u5_mult_82_ab_45__0_) );
  NOR2_X1 u5_mult_82_U1221 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n227), .ZN(
        u5_mult_82_ab_45__10_) );
  NOR2_X1 u5_mult_82_U1220 ( .A1(u5_mult_82_n426), .A2(u5_mult_82_n226), .ZN(
        u5_mult_82_ab_45__11_) );
  NOR2_X1 u5_mult_82_U1219 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n226), .ZN(
        u5_mult_82_ab_45__12_) );
  NOR2_X1 u5_mult_82_U1218 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n228), .ZN(
        u5_mult_82_ab_45__13_) );
  NOR2_X1 u5_mult_82_U1217 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n452), .ZN(
        u5_mult_82_ab_45__14_) );
  NOR2_X1 u5_mult_82_U1216 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n452), .ZN(
        u5_mult_82_ab_45__15_) );
  NOR2_X1 u5_mult_82_U1215 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n452), .ZN(
        u5_mult_82_ab_45__16_) );
  NOR2_X1 u5_mult_82_U1214 ( .A1(u5_mult_82_n409), .A2(u5_mult_82_n452), .ZN(
        u5_mult_82_ab_45__17_) );
  NOR2_X1 u5_mult_82_U1213 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n452), .ZN(
        u5_mult_82_ab_45__18_) );
  NOR2_X1 u5_mult_82_U1212 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n452), .ZN(
        u5_mult_82_ab_45__19_) );
  NOR2_X1 u5_mult_82_U1211 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n226), .ZN(
        u5_mult_82_ab_45__1_) );
  NOR2_X1 u5_mult_82_U1210 ( .A1(u5_mult_82_n475), .A2(u5_mult_82_n226), .ZN(
        u5_mult_82_ab_45__20_) );
  NOR2_X1 u5_mult_82_U1209 ( .A1(u5_mult_82_n402), .A2(u5_mult_82_n226), .ZN(
        u5_mult_82_ab_45__21_) );
  NOR2_X1 u5_mult_82_U1208 ( .A1(u5_mult_82_n400), .A2(u5_mult_82_n226), .ZN(
        u5_mult_82_ab_45__22_) );
  NOR2_X1 u5_mult_82_U1207 ( .A1(u5_mult_82_n398), .A2(u5_mult_82_n226), .ZN(
        u5_mult_82_ab_45__23_) );
  NOR2_X1 u5_mult_82_U1206 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n226), .ZN(
        u5_mult_82_ab_45__24_) );
  NOR2_X1 u5_mult_82_U1205 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n226), .ZN(
        u5_mult_82_ab_45__25_) );
  NOR2_X1 u5_mult_82_U1204 ( .A1(u5_mult_82_n392), .A2(u5_mult_82_n226), .ZN(
        u5_mult_82_ab_45__26_) );
  NOR2_X1 u5_mult_82_U1203 ( .A1(u5_mult_82_n390), .A2(u5_mult_82_n226), .ZN(
        u5_mult_82_ab_45__27_) );
  NOR2_X1 u5_mult_82_U1202 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n226), .ZN(
        u5_mult_82_ab_45__28_) );
  NOR2_X1 u5_mult_82_U1201 ( .A1(u5_mult_82_n386), .A2(u5_mult_82_n226), .ZN(
        u5_mult_82_ab_45__29_) );
  NOR2_X1 u5_mult_82_U1200 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n227), .ZN(
        u5_mult_82_ab_45__2_) );
  NOR2_X1 u5_mult_82_U1199 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n227), .ZN(
        u5_mult_82_ab_45__30_) );
  NOR2_X1 u5_mult_82_U1198 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n227), .ZN(
        u5_mult_82_ab_45__31_) );
  NOR2_X1 u5_mult_82_U1197 ( .A1(u5_mult_82_n380), .A2(u5_mult_82_n227), .ZN(
        u5_mult_82_ab_45__32_) );
  NOR2_X1 u5_mult_82_U1196 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n227), .ZN(
        u5_mult_82_ab_45__33_) );
  NOR2_X1 u5_mult_82_U1195 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n227), .ZN(
        u5_mult_82_ab_45__34_) );
  NOR2_X1 u5_mult_82_U1194 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n227), .ZN(
        u5_mult_82_ab_45__35_) );
  NOR2_X1 u5_mult_82_U1193 ( .A1(u5_mult_82_n474), .A2(u5_mult_82_n227), .ZN(
        u5_mult_82_ab_45__36_) );
  NOR2_X1 u5_mult_82_U1192 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n227), .ZN(
        u5_mult_82_ab_45__37_) );
  NOR2_X1 u5_mult_82_U1191 ( .A1(u5_mult_82_n367), .A2(u5_mult_82_n227), .ZN(
        u5_mult_82_ab_45__38_) );
  NOR2_X1 u5_mult_82_U1190 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n227), .ZN(
        u5_mult_82_ab_45__39_) );
  NOR2_X1 u5_mult_82_U1189 ( .A1(u5_mult_82_n478), .A2(u5_mult_82_n228), .ZN(
        u5_mult_82_ab_45__3_) );
  NOR2_X1 u5_mult_82_U1188 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n228), .ZN(
        u5_mult_82_ab_45__40_) );
  NOR2_X1 u5_mult_82_U1187 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n228), .ZN(
        u5_mult_82_ab_45__41_) );
  NOR2_X1 u5_mult_82_U1186 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n228), .ZN(
        u5_mult_82_ab_45__42_) );
  NOR2_X1 u5_mult_82_U1185 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n228), .ZN(
        u5_mult_82_ab_45__43_) );
  NOR2_X1 u5_mult_82_U1184 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n228), .ZN(
        u5_mult_82_ab_45__44_) );
  NOR2_X1 u5_mult_82_U1183 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n228), .ZN(
        u5_mult_82_ab_45__45_) );
  NOR2_X1 u5_mult_82_U1182 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n228), .ZN(
        u5_mult_82_ab_45__46_) );
  NOR2_X1 u5_mult_82_U1181 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n228), .ZN(
        u5_mult_82_ab_45__47_) );
  NOR2_X1 u5_mult_82_U1180 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n228), .ZN(
        u5_mult_82_ab_45__48_) );
  NOR2_X1 u5_mult_82_U1179 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n228), .ZN(
        u5_mult_82_ab_45__49_) );
  NOR2_X1 u5_mult_82_U1178 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n226), .ZN(
        u5_mult_82_ab_45__4_) );
  NOR2_X1 u5_mult_82_U1177 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n226), .ZN(
        u5_mult_82_ab_45__50_) );
  NOR2_X1 u5_mult_82_U1176 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n226), .ZN(
        u5_mult_82_ab_45__51_) );
  NOR2_X1 u5_mult_82_U1175 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n226), .ZN(
        u5_mult_82_ab_45__52_) );
  NOR2_X1 u5_mult_82_U1174 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n226), .ZN(
        u5_mult_82_ab_45__5_) );
  NOR2_X1 u5_mult_82_U1173 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n226), .ZN(
        u5_mult_82_ab_45__6_) );
  NOR2_X1 u5_mult_82_U1172 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n226), .ZN(
        u5_mult_82_ab_45__7_) );
  NOR2_X1 u5_mult_82_U1171 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n227), .ZN(
        u5_mult_82_ab_45__8_) );
  NOR2_X1 u5_mult_82_U1170 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n228), .ZN(
        u5_mult_82_ab_45__9_) );
  NOR2_X1 u5_mult_82_U1169 ( .A1(u5_mult_82_n480), .A2(u5_mult_82_n224), .ZN(
        u5_mult_82_ab_46__0_) );
  NOR2_X1 u5_mult_82_U1168 ( .A1(u5_mult_82_n477), .A2(u5_mult_82_n224), .ZN(
        u5_mult_82_ab_46__10_) );
  NOR2_X1 u5_mult_82_U1167 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n224), .ZN(
        u5_mult_82_ab_46__11_) );
  NOR2_X1 u5_mult_82_U1166 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n224), .ZN(
        u5_mult_82_ab_46__12_) );
  NOR2_X1 u5_mult_82_U1165 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n224), .ZN(
        u5_mult_82_ab_46__13_) );
  NOR2_X1 u5_mult_82_U1164 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n224), .ZN(
        u5_mult_82_ab_46__14_) );
  NOR2_X1 u5_mult_82_U1163 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n224), .ZN(
        u5_mult_82_ab_46__15_) );
  NOR2_X1 u5_mult_82_U1162 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n224), .ZN(
        u5_mult_82_ab_46__16_) );
  NOR2_X1 u5_mult_82_U1161 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n224), .ZN(
        u5_mult_82_ab_46__17_) );
  NOR2_X1 u5_mult_82_U1160 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n224), .ZN(
        u5_mult_82_ab_46__18_) );
  NOR2_X1 u5_mult_82_U1159 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n224), .ZN(
        u5_mult_82_ab_46__19_) );
  NOR2_X1 u5_mult_82_U1158 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n225), .ZN(
        u5_mult_82_ab_46__1_) );
  NOR2_X1 u5_mult_82_U1157 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n225), .ZN(
        u5_mult_82_ab_46__20_) );
  NOR2_X1 u5_mult_82_U1156 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n225), .ZN(
        u5_mult_82_ab_46__21_) );
  NOR2_X1 u5_mult_82_U1155 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n225), .ZN(
        u5_mult_82_ab_46__22_) );
  NOR2_X1 u5_mult_82_U1154 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n225), .ZN(
        u5_mult_82_ab_46__23_) );
  NOR2_X1 u5_mult_82_U1153 ( .A1(u5_mult_82_n396), .A2(u5_mult_82_n225), .ZN(
        u5_mult_82_ab_46__24_) );
  NOR2_X1 u5_mult_82_U1152 ( .A1(u5_mult_82_n394), .A2(u5_mult_82_n225), .ZN(
        u5_mult_82_ab_46__25_) );
  NOR2_X1 u5_mult_82_U1151 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n225), .ZN(
        u5_mult_82_ab_46__26_) );
  NOR2_X1 u5_mult_82_U1150 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n225), .ZN(
        u5_mult_82_ab_46__27_) );
  NOR2_X1 u5_mult_82_U1149 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n225), .ZN(
        u5_mult_82_ab_46__28_) );
  NOR2_X1 u5_mult_82_U1148 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n225), .ZN(
        u5_mult_82_ab_46__29_) );
  NOR2_X1 u5_mult_82_U1147 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n225), .ZN(
        u5_mult_82_ab_46__2_) );
  NOR2_X1 u5_mult_82_U1146 ( .A1(u5_mult_82_n384), .A2(u5_mult_82_n225), .ZN(
        u5_mult_82_ab_46__30_) );
  NOR2_X1 u5_mult_82_U1145 ( .A1(u5_mult_82_n382), .A2(u5_mult_82_n225), .ZN(
        u5_mult_82_ab_46__31_) );
  NOR2_X1 u5_mult_82_U1144 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n225), .ZN(
        u5_mult_82_ab_46__32_) );
  NOR2_X1 u5_mult_82_U1143 ( .A1(u5_mult_82_n378), .A2(u5_mult_82_n225), .ZN(
        u5_mult_82_ab_46__33_) );
  NOR2_X1 u5_mult_82_U1142 ( .A1(u5_mult_82_n376), .A2(u5_mult_82_n225), .ZN(
        u5_mult_82_ab_46__34_) );
  NOR2_X1 u5_mult_82_U1141 ( .A1(u5_mult_82_n374), .A2(u5_mult_82_n225), .ZN(
        u5_mult_82_ab_46__35_) );
  NOR2_X1 u5_mult_82_U1140 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n225), .ZN(
        u5_mult_82_ab_46__36_) );
  NOR2_X1 u5_mult_82_U1139 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n225), .ZN(
        u5_mult_82_ab_46__37_) );
  NOR2_X1 u5_mult_82_U1138 ( .A1(u5_mult_82_n367), .A2(u5_mult_82_n225), .ZN(
        u5_mult_82_ab_46__38_) );
  NOR2_X1 u5_mult_82_U1137 ( .A1(u5_mult_82_n366), .A2(u5_mult_82_n225), .ZN(
        u5_mult_82_ab_46__39_) );
  NOR2_X1 u5_mult_82_U1136 ( .A1(u5_mult_82_n478), .A2(u5_mult_82_n224), .ZN(
        u5_mult_82_ab_46__3_) );
  NOR2_X1 u5_mult_82_U1135 ( .A1(u5_mult_82_n364), .A2(u5_mult_82_n224), .ZN(
        u5_mult_82_ab_46__40_) );
  NOR2_X1 u5_mult_82_U1134 ( .A1(u5_mult_82_n362), .A2(u5_mult_82_n224), .ZN(
        u5_mult_82_ab_46__41_) );
  NOR2_X1 u5_mult_82_U1133 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n224), .ZN(
        u5_mult_82_ab_46__42_) );
  NOR2_X1 u5_mult_82_U1132 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n224), .ZN(
        u5_mult_82_ab_46__43_) );
  NOR2_X1 u5_mult_82_U1131 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n224), .ZN(
        u5_mult_82_ab_46__44_) );
  NOR2_X1 u5_mult_82_U1130 ( .A1(u5_mult_82_n352), .A2(u5_mult_82_n224), .ZN(
        u5_mult_82_ab_46__45_) );
  NOR2_X1 u5_mult_82_U1129 ( .A1(u5_mult_82_n350), .A2(u5_mult_82_n224), .ZN(
        u5_mult_82_ab_46__46_) );
  NOR2_X1 u5_mult_82_U1128 ( .A1(u5_mult_82_n348), .A2(u5_mult_82_n224), .ZN(
        u5_mult_82_ab_46__47_) );
  NOR2_X1 u5_mult_82_U1127 ( .A1(u5_mult_82_n346), .A2(u5_mult_82_n224), .ZN(
        u5_mult_82_ab_46__48_) );
  NOR2_X1 u5_mult_82_U1126 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n224), .ZN(
        u5_mult_82_ab_46__49_) );
  NOR2_X1 u5_mult_82_U1125 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n225), .ZN(
        u5_mult_82_ab_46__4_) );
  NOR2_X1 u5_mult_82_U1124 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n225), .ZN(
        u5_mult_82_ab_46__50_) );
  NOR2_X1 u5_mult_82_U1123 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n225), .ZN(
        u5_mult_82_ab_46__51_) );
  NOR2_X1 u5_mult_82_U1122 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n451), .ZN(
        u5_mult_82_ab_46__52_) );
  NOR2_X1 u5_mult_82_U1121 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n225), .ZN(
        u5_mult_82_ab_46__5_) );
  NOR2_X1 u5_mult_82_U1120 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n451), .ZN(
        u5_mult_82_ab_46__6_) );
  NOR2_X1 u5_mult_82_U1119 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n451), .ZN(
        u5_mult_82_ab_46__7_) );
  NOR2_X1 u5_mult_82_U1118 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n451), .ZN(
        u5_mult_82_ab_46__8_) );
  NOR2_X1 u5_mult_82_U1117 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n451), .ZN(
        u5_mult_82_ab_46__9_) );
  NOR2_X1 u5_mult_82_U1116 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n221), .ZN(
        u5_mult_82_ab_47__0_) );
  NOR2_X1 u5_mult_82_U1115 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n221), .ZN(
        u5_mult_82_ab_47__10_) );
  NOR2_X1 u5_mult_82_U1114 ( .A1(u5_mult_82_n426), .A2(u5_mult_82_n221), .ZN(
        u5_mult_82_ab_47__11_) );
  NOR2_X1 u5_mult_82_U1113 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n221), .ZN(
        u5_mult_82_ab_47__12_) );
  NOR2_X1 u5_mult_82_U1112 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n221), .ZN(
        u5_mult_82_ab_47__13_) );
  NOR2_X1 u5_mult_82_U1111 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n221), .ZN(
        u5_mult_82_ab_47__14_) );
  NOR2_X1 u5_mult_82_U1110 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n221), .ZN(
        u5_mult_82_ab_47__15_) );
  NOR2_X1 u5_mult_82_U1109 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n221), .ZN(
        u5_mult_82_ab_47__16_) );
  NOR2_X1 u5_mult_82_U1108 ( .A1(u5_mult_82_n409), .A2(u5_mult_82_n221), .ZN(
        u5_mult_82_ab_47__17_) );
  NOR2_X1 u5_mult_82_U1107 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n221), .ZN(
        u5_mult_82_ab_47__18_) );
  NOR2_X1 u5_mult_82_U1106 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n221), .ZN(
        u5_mult_82_ab_47__19_) );
  NOR2_X1 u5_mult_82_U1105 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n221), .ZN(
        u5_mult_82_ab_47__1_) );
  NOR2_X1 u5_mult_82_U1104 ( .A1(u5_mult_82_n475), .A2(u5_mult_82_n221), .ZN(
        u5_mult_82_ab_47__20_) );
  NOR2_X1 u5_mult_82_U1103 ( .A1(u5_mult_82_n402), .A2(u5_mult_82_n221), .ZN(
        u5_mult_82_ab_47__21_) );
  NOR2_X1 u5_mult_82_U1102 ( .A1(u5_mult_82_n400), .A2(u5_mult_82_n221), .ZN(
        u5_mult_82_ab_47__22_) );
  NOR2_X1 u5_mult_82_U1101 ( .A1(u5_mult_82_n398), .A2(u5_mult_82_n221), .ZN(
        u5_mult_82_ab_47__23_) );
  NOR2_X1 u5_mult_82_U1100 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n221), .ZN(
        u5_mult_82_ab_47__24_) );
  NOR2_X1 u5_mult_82_U1099 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n221), .ZN(
        u5_mult_82_ab_47__25_) );
  NOR2_X1 u5_mult_82_U1098 ( .A1(u5_mult_82_n392), .A2(u5_mult_82_n221), .ZN(
        u5_mult_82_ab_47__26_) );
  NOR2_X1 u5_mult_82_U1097 ( .A1(u5_mult_82_n390), .A2(u5_mult_82_n221), .ZN(
        u5_mult_82_ab_47__27_) );
  NOR2_X1 u5_mult_82_U1096 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n221), .ZN(
        u5_mult_82_ab_47__28_) );
  NOR2_X1 u5_mult_82_U1095 ( .A1(u5_mult_82_n386), .A2(u5_mult_82_n221), .ZN(
        u5_mult_82_ab_47__29_) );
  NOR2_X1 u5_mult_82_U1094 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n222), .ZN(
        u5_mult_82_ab_47__2_) );
  NOR2_X1 u5_mult_82_U1093 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n222), .ZN(
        u5_mult_82_ab_47__30_) );
  NOR2_X1 u5_mult_82_U1092 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n222), .ZN(
        u5_mult_82_ab_47__31_) );
  NOR2_X1 u5_mult_82_U1091 ( .A1(u5_mult_82_n380), .A2(u5_mult_82_n222), .ZN(
        u5_mult_82_ab_47__32_) );
  NOR2_X1 u5_mult_82_U1090 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n222), .ZN(
        u5_mult_82_ab_47__33_) );
  NOR2_X1 u5_mult_82_U1089 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n222), .ZN(
        u5_mult_82_ab_47__34_) );
  NOR2_X1 u5_mult_82_U1088 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n222), .ZN(
        u5_mult_82_ab_47__35_) );
  NOR2_X1 u5_mult_82_U1087 ( .A1(u5_mult_82_n474), .A2(u5_mult_82_n222), .ZN(
        u5_mult_82_ab_47__36_) );
  NOR2_X1 u5_mult_82_U1086 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n222), .ZN(
        u5_mult_82_ab_47__37_) );
  NOR2_X1 u5_mult_82_U1085 ( .A1(u5_mult_82_n367), .A2(u5_mult_82_n222), .ZN(
        u5_mult_82_ab_47__38_) );
  NOR2_X1 u5_mult_82_U1084 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n222), .ZN(
        u5_mult_82_ab_47__39_) );
  NOR2_X1 u5_mult_82_U1083 ( .A1(u5_mult_82_n478), .A2(u5_mult_82_n223), .ZN(
        u5_mult_82_ab_47__3_) );
  NOR2_X1 u5_mult_82_U1082 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n223), .ZN(
        u5_mult_82_ab_47__40_) );
  NOR2_X1 u5_mult_82_U1081 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n223), .ZN(
        u5_mult_82_ab_47__41_) );
  NOR2_X1 u5_mult_82_U1080 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n223), .ZN(
        u5_mult_82_ab_47__42_) );
  NOR2_X1 u5_mult_82_U1079 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n223), .ZN(
        u5_mult_82_ab_47__43_) );
  NOR2_X1 u5_mult_82_U1078 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n223), .ZN(
        u5_mult_82_ab_47__44_) );
  NOR2_X1 u5_mult_82_U1077 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n223), .ZN(
        u5_mult_82_ab_47__45_) );
  NOR2_X1 u5_mult_82_U1076 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n223), .ZN(
        u5_mult_82_ab_47__46_) );
  NOR2_X1 u5_mult_82_U1075 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n223), .ZN(
        u5_mult_82_ab_47__47_) );
  NOR2_X1 u5_mult_82_U1074 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n223), .ZN(
        u5_mult_82_ab_47__48_) );
  NOR2_X1 u5_mult_82_U1073 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n223), .ZN(
        u5_mult_82_ab_47__49_) );
  NOR2_X1 u5_mult_82_U1072 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n221), .ZN(
        u5_mult_82_ab_47__4_) );
  NOR2_X1 u5_mult_82_U1071 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n221), .ZN(
        u5_mult_82_ab_47__50_) );
  NOR2_X1 u5_mult_82_U1070 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n221), .ZN(
        u5_mult_82_ab_47__51_) );
  NOR2_X1 u5_mult_82_U1069 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n221), .ZN(
        u5_mult_82_ab_47__52_) );
  NOR2_X1 u5_mult_82_U1068 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n222), .ZN(
        u5_mult_82_ab_47__5_) );
  NOR2_X1 u5_mult_82_U1067 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n223), .ZN(
        u5_mult_82_ab_47__6_) );
  NOR2_X1 u5_mult_82_U1066 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n222), .ZN(
        u5_mult_82_ab_47__7_) );
  NOR2_X1 u5_mult_82_U1065 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n222), .ZN(
        u5_mult_82_ab_47__8_) );
  NOR2_X1 u5_mult_82_U1064 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n221), .ZN(
        u5_mult_82_ab_47__9_) );
  NOR2_X1 u5_mult_82_U1063 ( .A1(u5_mult_82_n480), .A2(u5_mult_82_n218), .ZN(
        u5_mult_82_ab_48__0_) );
  NOR2_X1 u5_mult_82_U1062 ( .A1(u5_mult_82_n477), .A2(u5_mult_82_n218), .ZN(
        u5_mult_82_ab_48__10_) );
  NOR2_X1 u5_mult_82_U1061 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n218), .ZN(
        u5_mult_82_ab_48__11_) );
  NOR2_X1 u5_mult_82_U1060 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n218), .ZN(
        u5_mult_82_ab_48__12_) );
  NOR2_X1 u5_mult_82_U1059 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n218), .ZN(
        u5_mult_82_ab_48__13_) );
  NOR2_X1 u5_mult_82_U1058 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n218), .ZN(
        u5_mult_82_ab_48__14_) );
  NOR2_X1 u5_mult_82_U1057 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n218), .ZN(
        u5_mult_82_ab_48__15_) );
  NOR2_X1 u5_mult_82_U1056 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n218), .ZN(
        u5_mult_82_ab_48__16_) );
  NOR2_X1 u5_mult_82_U1055 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n218), .ZN(
        u5_mult_82_ab_48__17_) );
  NOR2_X1 u5_mult_82_U1054 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n218), .ZN(
        u5_mult_82_ab_48__18_) );
  NOR2_X1 u5_mult_82_U1053 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n218), .ZN(
        u5_mult_82_ab_48__19_) );
  NOR2_X1 u5_mult_82_U1052 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n218), .ZN(
        u5_mult_82_ab_48__1_) );
  NOR2_X1 u5_mult_82_U1051 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n218), .ZN(
        u5_mult_82_ab_48__20_) );
  NOR2_X1 u5_mult_82_U1050 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n218), .ZN(
        u5_mult_82_ab_48__21_) );
  NOR2_X1 u5_mult_82_U1049 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n218), .ZN(
        u5_mult_82_ab_48__22_) );
  NOR2_X1 u5_mult_82_U1048 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n218), .ZN(
        u5_mult_82_ab_48__23_) );
  NOR2_X1 u5_mult_82_U1047 ( .A1(u5_mult_82_n396), .A2(u5_mult_82_n218), .ZN(
        u5_mult_82_ab_48__24_) );
  NOR2_X1 u5_mult_82_U1046 ( .A1(u5_mult_82_n394), .A2(u5_mult_82_n218), .ZN(
        u5_mult_82_ab_48__25_) );
  NOR2_X1 u5_mult_82_U1045 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n218), .ZN(
        u5_mult_82_ab_48__26_) );
  NOR2_X1 u5_mult_82_U1044 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n218), .ZN(
        u5_mult_82_ab_48__27_) );
  NOR2_X1 u5_mult_82_U1043 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n218), .ZN(
        u5_mult_82_ab_48__28_) );
  NOR2_X1 u5_mult_82_U1042 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n218), .ZN(
        u5_mult_82_ab_48__29_) );
  NOR2_X1 u5_mult_82_U1041 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n219), .ZN(
        u5_mult_82_ab_48__2_) );
  NOR2_X1 u5_mult_82_U1040 ( .A1(u5_mult_82_n384), .A2(u5_mult_82_n219), .ZN(
        u5_mult_82_ab_48__30_) );
  NOR2_X1 u5_mult_82_U1039 ( .A1(u5_mult_82_n382), .A2(u5_mult_82_n219), .ZN(
        u5_mult_82_ab_48__31_) );
  NOR2_X1 u5_mult_82_U1038 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n219), .ZN(
        u5_mult_82_ab_48__32_) );
  NOR2_X1 u5_mult_82_U1037 ( .A1(u5_mult_82_n378), .A2(u5_mult_82_n219), .ZN(
        u5_mult_82_ab_48__33_) );
  NOR2_X1 u5_mult_82_U1036 ( .A1(u5_mult_82_n376), .A2(u5_mult_82_n219), .ZN(
        u5_mult_82_ab_48__34_) );
  NOR2_X1 u5_mult_82_U1035 ( .A1(u5_mult_82_n374), .A2(u5_mult_82_n219), .ZN(
        u5_mult_82_ab_48__35_) );
  NOR2_X1 u5_mult_82_U1034 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n219), .ZN(
        u5_mult_82_ab_48__36_) );
  NOR2_X1 u5_mult_82_U1033 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n219), .ZN(
        u5_mult_82_ab_48__37_) );
  NOR2_X1 u5_mult_82_U1032 ( .A1(u5_mult_82_n367), .A2(u5_mult_82_n219), .ZN(
        u5_mult_82_ab_48__38_) );
  NOR2_X1 u5_mult_82_U1031 ( .A1(u5_mult_82_n366), .A2(u5_mult_82_n219), .ZN(
        u5_mult_82_ab_48__39_) );
  NOR2_X1 u5_mult_82_U1030 ( .A1(u5_mult_82_n478), .A2(u5_mult_82_n220), .ZN(
        u5_mult_82_ab_48__3_) );
  NOR2_X1 u5_mult_82_U1029 ( .A1(u5_mult_82_n364), .A2(u5_mult_82_n220), .ZN(
        u5_mult_82_ab_48__40_) );
  NOR2_X1 u5_mult_82_U1028 ( .A1(u5_mult_82_n362), .A2(u5_mult_82_n220), .ZN(
        u5_mult_82_ab_48__41_) );
  NOR2_X1 u5_mult_82_U1027 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n220), .ZN(
        u5_mult_82_ab_48__42_) );
  NOR2_X1 u5_mult_82_U1026 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n220), .ZN(
        u5_mult_82_ab_48__43_) );
  NOR2_X1 u5_mult_82_U1025 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n220), .ZN(
        u5_mult_82_ab_48__44_) );
  NOR2_X1 u5_mult_82_U1024 ( .A1(u5_mult_82_n352), .A2(u5_mult_82_n220), .ZN(
        u5_mult_82_ab_48__45_) );
  NOR2_X1 u5_mult_82_U1023 ( .A1(u5_mult_82_n350), .A2(u5_mult_82_n220), .ZN(
        u5_mult_82_ab_48__46_) );
  NOR2_X1 u5_mult_82_U1022 ( .A1(u5_mult_82_n348), .A2(u5_mult_82_n220), .ZN(
        u5_mult_82_ab_48__47_) );
  NOR2_X1 u5_mult_82_U1021 ( .A1(u5_mult_82_n346), .A2(u5_mult_82_n220), .ZN(
        u5_mult_82_ab_48__48_) );
  NOR2_X1 u5_mult_82_U1020 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n220), .ZN(
        u5_mult_82_ab_48__49_) );
  NOR2_X1 u5_mult_82_U1019 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n220), .ZN(
        u5_mult_82_ab_48__4_) );
  NOR2_X1 u5_mult_82_U1018 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n218), .ZN(
        u5_mult_82_ab_48__50_) );
  NOR2_X1 u5_mult_82_U1017 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n218), .ZN(
        u5_mult_82_ab_48__51_) );
  NOR2_X1 u5_mult_82_U1016 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n218), .ZN(
        u5_mult_82_ab_48__52_) );
  NOR2_X1 u5_mult_82_U1015 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n219), .ZN(
        u5_mult_82_ab_48__5_) );
  NOR2_X1 u5_mult_82_U1014 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n220), .ZN(
        u5_mult_82_ab_48__6_) );
  NOR2_X1 u5_mult_82_U1013 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n219), .ZN(
        u5_mult_82_ab_48__7_) );
  NOR2_X1 u5_mult_82_U1012 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n219), .ZN(
        u5_mult_82_ab_48__8_) );
  NOR2_X1 u5_mult_82_U1011 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n218), .ZN(
        u5_mult_82_ab_48__9_) );
  NOR2_X1 u5_mult_82_U1010 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n215), .ZN(
        u5_mult_82_ab_49__0_) );
  NOR2_X1 u5_mult_82_U1009 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n215), .ZN(
        u5_mult_82_ab_49__10_) );
  NOR2_X1 u5_mult_82_U1008 ( .A1(u5_mult_82_n426), .A2(u5_mult_82_n215), .ZN(
        u5_mult_82_ab_49__11_) );
  NOR2_X1 u5_mult_82_U1007 ( .A1(u5_mult_82_n423), .A2(u5_mult_82_n215), .ZN(
        u5_mult_82_ab_49__12_) );
  NOR2_X1 u5_mult_82_U1006 ( .A1(u5_mult_82_n420), .A2(u5_mult_82_n215), .ZN(
        u5_mult_82_ab_49__13_) );
  NOR2_X1 u5_mult_82_U1005 ( .A1(u5_mult_82_n417), .A2(u5_mult_82_n215), .ZN(
        u5_mult_82_ab_49__14_) );
  NOR2_X1 u5_mult_82_U1004 ( .A1(u5_mult_82_n414), .A2(u5_mult_82_n215), .ZN(
        u5_mult_82_ab_49__15_) );
  NOR2_X1 u5_mult_82_U1003 ( .A1(u5_mult_82_n411), .A2(u5_mult_82_n215), .ZN(
        u5_mult_82_ab_49__16_) );
  NOR2_X1 u5_mult_82_U1002 ( .A1(u5_mult_82_n409), .A2(u5_mult_82_n215), .ZN(
        u5_mult_82_ab_49__17_) );
  NOR2_X1 u5_mult_82_U1001 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n215), .ZN(
        u5_mult_82_ab_49__18_) );
  NOR2_X1 u5_mult_82_U1000 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n215), .ZN(
        u5_mult_82_ab_49__19_) );
  NOR2_X1 u5_mult_82_U999 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n215), .ZN(
        u5_mult_82_ab_49__1_) );
  NOR2_X1 u5_mult_82_U998 ( .A1(u5_mult_82_n475), .A2(u5_mult_82_n215), .ZN(
        u5_mult_82_ab_49__20_) );
  NOR2_X1 u5_mult_82_U997 ( .A1(u5_mult_82_n402), .A2(u5_mult_82_n215), .ZN(
        u5_mult_82_ab_49__21_) );
  NOR2_X1 u5_mult_82_U996 ( .A1(u5_mult_82_n400), .A2(u5_mult_82_n215), .ZN(
        u5_mult_82_ab_49__22_) );
  NOR2_X1 u5_mult_82_U995 ( .A1(u5_mult_82_n398), .A2(u5_mult_82_n215), .ZN(
        u5_mult_82_ab_49__23_) );
  NOR2_X1 u5_mult_82_U994 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n215), .ZN(
        u5_mult_82_ab_49__24_) );
  NOR2_X1 u5_mult_82_U993 ( .A1(u5_mult_82_n394), .A2(u5_mult_82_n215), .ZN(
        u5_mult_82_ab_49__25_) );
  NOR2_X1 u5_mult_82_U992 ( .A1(u5_mult_82_n392), .A2(u5_mult_82_n215), .ZN(
        u5_mult_82_ab_49__26_) );
  NOR2_X1 u5_mult_82_U991 ( .A1(u5_mult_82_n390), .A2(u5_mult_82_n215), .ZN(
        u5_mult_82_ab_49__27_) );
  NOR2_X1 u5_mult_82_U990 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n215), .ZN(
        u5_mult_82_ab_49__28_) );
  NOR2_X1 u5_mult_82_U989 ( .A1(u5_mult_82_n386), .A2(u5_mult_82_n215), .ZN(
        u5_mult_82_ab_49__29_) );
  NOR2_X1 u5_mult_82_U988 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n216), .ZN(
        u5_mult_82_ab_49__2_) );
  NOR2_X1 u5_mult_82_U987 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n216), .ZN(
        u5_mult_82_ab_49__30_) );
  NOR2_X1 u5_mult_82_U986 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n216), .ZN(
        u5_mult_82_ab_49__31_) );
  NOR2_X1 u5_mult_82_U985 ( .A1(u5_mult_82_n380), .A2(u5_mult_82_n216), .ZN(
        u5_mult_82_ab_49__32_) );
  NOR2_X1 u5_mult_82_U984 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n216), .ZN(
        u5_mult_82_ab_49__33_) );
  NOR2_X1 u5_mult_82_U983 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n216), .ZN(
        u5_mult_82_ab_49__34_) );
  NOR2_X1 u5_mult_82_U982 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n216), .ZN(
        u5_mult_82_ab_49__35_) );
  NOR2_X1 u5_mult_82_U981 ( .A1(u5_mult_82_n474), .A2(u5_mult_82_n216), .ZN(
        u5_mult_82_ab_49__36_) );
  NOR2_X1 u5_mult_82_U980 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n216), .ZN(
        u5_mult_82_ab_49__37_) );
  NOR2_X1 u5_mult_82_U979 ( .A1(u5_mult_82_n367), .A2(u5_mult_82_n216), .ZN(
        u5_mult_82_ab_49__38_) );
  NOR2_X1 u5_mult_82_U978 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n216), .ZN(
        u5_mult_82_ab_49__39_) );
  NOR2_X1 u5_mult_82_U977 ( .A1(u5_mult_82_n478), .A2(u5_mult_82_n217), .ZN(
        u5_mult_82_ab_49__3_) );
  NOR2_X1 u5_mult_82_U976 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n217), .ZN(
        u5_mult_82_ab_49__40_) );
  NOR2_X1 u5_mult_82_U975 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n217), .ZN(
        u5_mult_82_ab_49__41_) );
  NOR2_X1 u5_mult_82_U974 ( .A1(u5_mult_82_n359), .A2(u5_mult_82_n217), .ZN(
        u5_mult_82_ab_49__42_) );
  NOR2_X1 u5_mult_82_U973 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n217), .ZN(
        u5_mult_82_ab_49__43_) );
  NOR2_X1 u5_mult_82_U972 ( .A1(u5_mult_82_n354), .A2(u5_mult_82_n217), .ZN(
        u5_mult_82_ab_49__44_) );
  NOR2_X1 u5_mult_82_U971 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n217), .ZN(
        u5_mult_82_ab_49__45_) );
  NOR2_X1 u5_mult_82_U970 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n217), .ZN(
        u5_mult_82_ab_49__46_) );
  NOR2_X1 u5_mult_82_U969 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n217), .ZN(
        u5_mult_82_ab_49__47_) );
  NOR2_X1 u5_mult_82_U968 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n217), .ZN(
        u5_mult_82_ab_49__48_) );
  NOR2_X1 u5_mult_82_U967 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n217), .ZN(
        u5_mult_82_ab_49__49_) );
  NOR2_X1 u5_mult_82_U966 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n217), .ZN(
        u5_mult_82_ab_49__4_) );
  NOR2_X1 u5_mult_82_U965 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n215), .ZN(
        u5_mult_82_ab_49__50_) );
  NOR2_X1 u5_mult_82_U964 ( .A1(u5_mult_82_n339), .A2(u5_mult_82_n215), .ZN(
        u5_mult_82_ab_49__51_) );
  NOR2_X1 u5_mult_82_U963 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n215), .ZN(
        u5_mult_82_ab_49__52_) );
  NOR2_X1 u5_mult_82_U962 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n216), .ZN(
        u5_mult_82_ab_49__5_) );
  NOR2_X1 u5_mult_82_U961 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n216), .ZN(
        u5_mult_82_ab_49__6_) );
  NOR2_X1 u5_mult_82_U960 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n216), .ZN(
        u5_mult_82_ab_49__7_) );
  NOR2_X1 u5_mult_82_U959 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n215), .ZN(
        u5_mult_82_ab_49__8_) );
  NOR2_X1 u5_mult_82_U958 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n215), .ZN(
        u5_mult_82_ab_49__9_) );
  NOR2_X1 u5_mult_82_U957 ( .A1(u5_mult_82_n480), .A2(u5_mult_82_n324), .ZN(
        u5_mult_82_ab_4__0_) );
  NOR2_X1 u5_mult_82_U956 ( .A1(u5_mult_82_n477), .A2(u5_mult_82_n324), .ZN(
        u5_mult_82_ab_4__10_) );
  NOR2_X1 u5_mult_82_U955 ( .A1(u5_mult_82_n426), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__11_) );
  NOR2_X1 u5_mult_82_U954 ( .A1(u5_mult_82_n424), .A2(u5_mult_82_n324), .ZN(
        u5_mult_82_ab_4__12_) );
  NOR2_X1 u5_mult_82_U953 ( .A1(u5_mult_82_n421), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__13_) );
  NOR2_X1 u5_mult_82_U952 ( .A1(u5_mult_82_n418), .A2(u5_mult_82_n324), .ZN(
        u5_mult_82_ab_4__14_) );
  NOR2_X1 u5_mult_82_U951 ( .A1(u5_mult_82_n415), .A2(u5_mult_82_n324), .ZN(
        u5_mult_82_ab_4__15_) );
  NOR2_X1 u5_mult_82_U950 ( .A1(u5_mult_82_n412), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__16_) );
  NOR2_X1 u5_mult_82_U949 ( .A1(u5_mult_82_n409), .A2(u5_mult_82_n324), .ZN(
        u5_mult_82_ab_4__17_) );
  NOR2_X1 u5_mult_82_U948 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__18_) );
  NOR2_X1 u5_mult_82_U947 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n324), .ZN(
        u5_mult_82_ab_4__19_) );
  NOR2_X1 u5_mult_82_U946 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__1_) );
  NOR2_X1 u5_mult_82_U945 ( .A1(u5_mult_82_n475), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__20_) );
  NOR2_X1 u5_mult_82_U944 ( .A1(u5_mult_82_n402), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__21_) );
  NOR2_X1 u5_mult_82_U943 ( .A1(u5_mult_82_n400), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__22_) );
  NOR2_X1 u5_mult_82_U942 ( .A1(u5_mult_82_n398), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__23_) );
  NOR2_X1 u5_mult_82_U941 ( .A1(u5_mult_82_n396), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__24_) );
  NOR2_X1 u5_mult_82_U940 ( .A1(u5_mult_82_n394), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__25_) );
  NOR2_X1 u5_mult_82_U939 ( .A1(u5_mult_82_n392), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__26_) );
  NOR2_X1 u5_mult_82_U938 ( .A1(u5_mult_82_n390), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__27_) );
  NOR2_X1 u5_mult_82_U937 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__28_) );
  NOR2_X1 u5_mult_82_U936 ( .A1(u5_mult_82_n386), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__29_) );
  NOR2_X1 u5_mult_82_U935 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__2_) );
  NOR2_X1 u5_mult_82_U934 ( .A1(u5_mult_82_n384), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__30_) );
  NOR2_X1 u5_mult_82_U933 ( .A1(u5_mult_82_n382), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__31_) );
  NOR2_X1 u5_mult_82_U932 ( .A1(u5_mult_82_n380), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__32_) );
  NOR2_X1 u5_mult_82_U931 ( .A1(u5_mult_82_n378), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__33_) );
  NOR2_X1 u5_mult_82_U930 ( .A1(u5_mult_82_n376), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__34_) );
  NOR2_X1 u5_mult_82_U929 ( .A1(u5_mult_82_n374), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__35_) );
  NOR2_X1 u5_mult_82_U928 ( .A1(u5_mult_82_n474), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__36_) );
  NOR2_X1 u5_mult_82_U927 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__37_) );
  NOR2_X1 u5_mult_82_U926 ( .A1(u5_mult_82_n368), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__38_) );
  NOR2_X1 u5_mult_82_U925 ( .A1(u5_mult_82_n366), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__39_) );
  NOR2_X1 u5_mult_82_U924 ( .A1(u5_mult_82_n441), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__3_) );
  NOR2_X1 u5_mult_82_U923 ( .A1(u5_mult_82_n364), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__40_) );
  NOR2_X1 u5_mult_82_U922 ( .A1(u5_mult_82_n362), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__41_) );
  NOR2_X1 u5_mult_82_U921 ( .A1(u5_mult_82_n360), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__42_) );
  NOR2_X1 u5_mult_82_U920 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__43_) );
  NOR2_X1 u5_mult_82_U919 ( .A1(u5_mult_82_n355), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__44_) );
  NOR2_X1 u5_mult_82_U918 ( .A1(u5_mult_82_n352), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__45_) );
  NOR2_X1 u5_mult_82_U917 ( .A1(u5_mult_82_n350), .A2(u5_mult_82_n324), .ZN(
        u5_mult_82_ab_4__46_) );
  NOR2_X1 u5_mult_82_U916 ( .A1(u5_mult_82_n348), .A2(u5_mult_82_n324), .ZN(
        u5_mult_82_ab_4__47_) );
  NOR2_X1 u5_mult_82_U915 ( .A1(u5_mult_82_n346), .A2(u5_mult_82_n324), .ZN(
        u5_mult_82_ab_4__48_) );
  NOR2_X1 u5_mult_82_U914 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n324), .ZN(
        u5_mult_82_ab_4__49_) );
  NOR2_X1 u5_mult_82_U913 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n324), .ZN(
        u5_mult_82_ab_4__4_) );
  NOR2_X1 u5_mult_82_U912 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n324), .ZN(
        u5_mult_82_ab_4__50_) );
  NOR2_X1 u5_mult_82_U911 ( .A1(u5_mult_82_n340), .A2(u5_mult_82_n324), .ZN(
        u5_mult_82_ab_4__51_) );
  NOR2_X1 u5_mult_82_U910 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__52_) );
  NOR2_X1 u5_mult_82_U909 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__5_) );
  NOR2_X1 u5_mult_82_U908 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n324), .ZN(
        u5_mult_82_ab_4__6_) );
  NOR2_X1 u5_mult_82_U907 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__7_) );
  NOR2_X1 u5_mult_82_U906 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n324), .ZN(
        u5_mult_82_ab_4__8_) );
  NOR2_X1 u5_mult_82_U905 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n323), .ZN(
        u5_mult_82_ab_4__9_) );
  NOR2_X1 u5_mult_82_U904 ( .A1(u5_mult_82_n480), .A2(u5_mult_82_n213), .ZN(
        u5_mult_82_ab_50__0_) );
  NOR2_X1 u5_mult_82_U903 ( .A1(u5_mult_82_n477), .A2(u5_mult_82_n213), .ZN(
        u5_mult_82_ab_50__10_) );
  NOR2_X1 u5_mult_82_U902 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n213), .ZN(
        u5_mult_82_ab_50__11_) );
  NOR2_X1 u5_mult_82_U901 ( .A1(u5_mult_82_n424), .A2(u5_mult_82_n213), .ZN(
        u5_mult_82_ab_50__12_) );
  NOR2_X1 u5_mult_82_U900 ( .A1(u5_mult_82_n421), .A2(u5_mult_82_n213), .ZN(
        u5_mult_82_ab_50__13_) );
  NOR2_X1 u5_mult_82_U899 ( .A1(u5_mult_82_n418), .A2(u5_mult_82_n213), .ZN(
        u5_mult_82_ab_50__14_) );
  NOR2_X1 u5_mult_82_U898 ( .A1(u5_mult_82_n415), .A2(u5_mult_82_n213), .ZN(
        u5_mult_82_ab_50__15_) );
  NOR2_X1 u5_mult_82_U897 ( .A1(u5_mult_82_n412), .A2(u5_mult_82_n213), .ZN(
        u5_mult_82_ab_50__16_) );
  NOR2_X1 u5_mult_82_U896 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n213), .ZN(
        u5_mult_82_ab_50__17_) );
  NOR2_X1 u5_mult_82_U895 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n213), .ZN(
        u5_mult_82_ab_50__18_) );
  NOR2_X1 u5_mult_82_U894 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n213), .ZN(
        u5_mult_82_ab_50__19_) );
  NOR2_X1 u5_mult_82_U893 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n213), .ZN(
        u5_mult_82_ab_50__1_) );
  NOR2_X1 u5_mult_82_U892 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n213), .ZN(
        u5_mult_82_ab_50__20_) );
  NOR2_X1 u5_mult_82_U891 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n213), .ZN(
        u5_mult_82_ab_50__21_) );
  NOR2_X1 u5_mult_82_U890 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n213), .ZN(
        u5_mult_82_ab_50__22_) );
  NOR2_X1 u5_mult_82_U889 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n213), .ZN(
        u5_mult_82_ab_50__23_) );
  NOR2_X1 u5_mult_82_U888 ( .A1(u5_mult_82_n396), .A2(u5_mult_82_n214), .ZN(
        u5_mult_82_ab_50__24_) );
  NOR2_X1 u5_mult_82_U887 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n213), .ZN(
        u5_mult_82_ab_50__25_) );
  NOR2_X1 u5_mult_82_U886 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n214), .ZN(
        u5_mult_82_ab_50__26_) );
  NOR2_X1 u5_mult_82_U885 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n214), .ZN(
        u5_mult_82_ab_50__27_) );
  NOR2_X1 u5_mult_82_U884 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n214), .ZN(
        u5_mult_82_ab_50__28_) );
  NOR2_X1 u5_mult_82_U883 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n450), .ZN(
        u5_mult_82_ab_50__29_) );
  NOR2_X1 u5_mult_82_U882 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n450), .ZN(
        u5_mult_82_ab_50__2_) );
  NOR2_X1 u5_mult_82_U881 ( .A1(u5_mult_82_n384), .A2(u5_mult_82_n450), .ZN(
        u5_mult_82_ab_50__30_) );
  NOR2_X1 u5_mult_82_U880 ( .A1(u5_mult_82_n382), .A2(u5_mult_82_n214), .ZN(
        u5_mult_82_ab_50__31_) );
  NOR2_X1 u5_mult_82_U879 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n450), .ZN(
        u5_mult_82_ab_50__32_) );
  NOR2_X1 u5_mult_82_U878 ( .A1(u5_mult_82_n378), .A2(u5_mult_82_n450), .ZN(
        u5_mult_82_ab_50__33_) );
  NOR2_X1 u5_mult_82_U877 ( .A1(u5_mult_82_n376), .A2(u5_mult_82_n450), .ZN(
        u5_mult_82_ab_50__34_) );
  NOR2_X1 u5_mult_82_U876 ( .A1(u5_mult_82_n374), .A2(u5_mult_82_n450), .ZN(
        u5_mult_82_ab_50__35_) );
  NOR2_X1 u5_mult_82_U875 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n213), .ZN(
        u5_mult_82_ab_50__36_) );
  NOR2_X1 u5_mult_82_U874 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n450), .ZN(
        u5_mult_82_ab_50__37_) );
  NOR2_X1 u5_mult_82_U873 ( .A1(u5_mult_82_n368), .A2(u5_mult_82_n214), .ZN(
        u5_mult_82_ab_50__38_) );
  NOR2_X1 u5_mult_82_U872 ( .A1(u5_mult_82_n366), .A2(u5_mult_82_n450), .ZN(
        u5_mult_82_ab_50__39_) );
  NOR2_X1 u5_mult_82_U871 ( .A1(u5_mult_82_n441), .A2(u5_mult_82_n214), .ZN(
        u5_mult_82_ab_50__3_) );
  NOR2_X1 u5_mult_82_U870 ( .A1(u5_mult_82_n364), .A2(u5_mult_82_n214), .ZN(
        u5_mult_82_ab_50__40_) );
  NOR2_X1 u5_mult_82_U869 ( .A1(u5_mult_82_n362), .A2(u5_mult_82_n214), .ZN(
        u5_mult_82_ab_50__41_) );
  NOR2_X1 u5_mult_82_U868 ( .A1(u5_mult_82_n360), .A2(u5_mult_82_n214), .ZN(
        u5_mult_82_ab_50__42_) );
  NOR2_X1 u5_mult_82_U867 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n214), .ZN(
        u5_mult_82_ab_50__43_) );
  NOR2_X1 u5_mult_82_U866 ( .A1(u5_mult_82_n355), .A2(u5_mult_82_n214), .ZN(
        u5_mult_82_ab_50__44_) );
  NOR2_X1 u5_mult_82_U865 ( .A1(u5_mult_82_n352), .A2(u5_mult_82_n214), .ZN(
        u5_mult_82_ab_50__45_) );
  NOR2_X1 u5_mult_82_U864 ( .A1(u5_mult_82_n350), .A2(u5_mult_82_n214), .ZN(
        u5_mult_82_ab_50__46_) );
  NOR2_X1 u5_mult_82_U863 ( .A1(u5_mult_82_n348), .A2(u5_mult_82_n214), .ZN(
        u5_mult_82_ab_50__47_) );
  NOR2_X1 u5_mult_82_U862 ( .A1(u5_mult_82_n346), .A2(u5_mult_82_n214), .ZN(
        u5_mult_82_ab_50__48_) );
  NOR2_X1 u5_mult_82_U861 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n214), .ZN(
        u5_mult_82_ab_50__49_) );
  NOR2_X1 u5_mult_82_U860 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n450), .ZN(
        u5_mult_82_ab_50__4_) );
  NOR2_X1 u5_mult_82_U859 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n213), .ZN(
        u5_mult_82_ab_50__50_) );
  NOR2_X1 u5_mult_82_U858 ( .A1(u5_mult_82_n340), .A2(u5_mult_82_n213), .ZN(
        u5_mult_82_ab_50__51_) );
  NOR2_X1 u5_mult_82_U857 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n213), .ZN(
        u5_mult_82_ab_50__52_) );
  NOR2_X1 u5_mult_82_U856 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n450), .ZN(
        u5_mult_82_ab_50__5_) );
  NOR2_X1 u5_mult_82_U855 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n213), .ZN(
        u5_mult_82_ab_50__6_) );
  NOR2_X1 u5_mult_82_U854 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n213), .ZN(
        u5_mult_82_ab_50__7_) );
  NOR2_X1 u5_mult_82_U853 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n213), .ZN(
        u5_mult_82_ab_50__8_) );
  NOR2_X1 u5_mult_82_U852 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n213), .ZN(
        u5_mult_82_ab_50__9_) );
  NOR2_X1 u5_mult_82_U851 ( .A1(u5_mult_82_n446), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__0_) );
  NOR2_X1 u5_mult_82_U850 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__10_) );
  NOR2_X1 u5_mult_82_U849 ( .A1(u5_mult_82_n426), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__11_) );
  NOR2_X1 u5_mult_82_U848 ( .A1(u5_mult_82_n424), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__12_) );
  NOR2_X1 u5_mult_82_U847 ( .A1(u5_mult_82_n421), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__13_) );
  NOR2_X1 u5_mult_82_U846 ( .A1(u5_mult_82_n418), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__14_) );
  NOR2_X1 u5_mult_82_U845 ( .A1(u5_mult_82_n415), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__15_) );
  NOR2_X1 u5_mult_82_U844 ( .A1(u5_mult_82_n412), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__16_) );
  NOR2_X1 u5_mult_82_U843 ( .A1(u5_mult_82_n409), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__17_) );
  NOR2_X1 u5_mult_82_U842 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__18_) );
  NOR2_X1 u5_mult_82_U841 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__19_) );
  NOR2_X1 u5_mult_82_U840 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n212), .ZN(
        u5_mult_82_ab_51__1_) );
  NOR2_X1 u5_mult_82_U839 ( .A1(u5_mult_82_n475), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__20_) );
  NOR2_X1 u5_mult_82_U838 ( .A1(u5_mult_82_n402), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__21_) );
  NOR2_X1 u5_mult_82_U837 ( .A1(u5_mult_82_n400), .A2(u5_mult_82_n212), .ZN(
        u5_mult_82_ab_51__22_) );
  NOR2_X1 u5_mult_82_U836 ( .A1(u5_mult_82_n398), .A2(u5_mult_82_n212), .ZN(
        u5_mult_82_ab_51__23_) );
  NOR2_X1 u5_mult_82_U835 ( .A1(u5_mult_82_n396), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__24_) );
  NOR2_X1 u5_mult_82_U834 ( .A1(u5_mult_82_n394), .A2(u5_mult_82_n212), .ZN(
        u5_mult_82_ab_51__25_) );
  NOR2_X1 u5_mult_82_U833 ( .A1(u5_mult_82_n392), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__26_) );
  NOR2_X1 u5_mult_82_U832 ( .A1(u5_mult_82_n390), .A2(u5_mult_82_n212), .ZN(
        u5_mult_82_ab_51__27_) );
  NOR2_X1 u5_mult_82_U831 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n212), .ZN(
        u5_mult_82_ab_51__28_) );
  NOR2_X1 u5_mult_82_U830 ( .A1(u5_mult_82_n386), .A2(u5_mult_82_n212), .ZN(
        u5_mult_82_ab_51__29_) );
  NOR2_X1 u5_mult_82_U829 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n212), .ZN(
        u5_mult_82_ab_51__2_) );
  NOR2_X1 u5_mult_82_U828 ( .A1(u5_mult_82_n383), .A2(u5_mult_82_n212), .ZN(
        u5_mult_82_ab_51__30_) );
  NOR2_X1 u5_mult_82_U827 ( .A1(u5_mult_82_n381), .A2(u5_mult_82_n212), .ZN(
        u5_mult_82_ab_51__31_) );
  NOR2_X1 u5_mult_82_U826 ( .A1(u5_mult_82_n380), .A2(u5_mult_82_n212), .ZN(
        u5_mult_82_ab_51__32_) );
  NOR2_X1 u5_mult_82_U825 ( .A1(u5_mult_82_n377), .A2(u5_mult_82_n212), .ZN(
        u5_mult_82_ab_51__33_) );
  NOR2_X1 u5_mult_82_U824 ( .A1(u5_mult_82_n375), .A2(u5_mult_82_n212), .ZN(
        u5_mult_82_ab_51__34_) );
  NOR2_X1 u5_mult_82_U823 ( .A1(u5_mult_82_n373), .A2(u5_mult_82_n212), .ZN(
        u5_mult_82_ab_51__35_) );
  NOR2_X1 u5_mult_82_U822 ( .A1(u5_mult_82_n474), .A2(u5_mult_82_n212), .ZN(
        u5_mult_82_ab_51__36_) );
  NOR2_X1 u5_mult_82_U821 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n212), .ZN(
        u5_mult_82_ab_51__37_) );
  NOR2_X1 u5_mult_82_U820 ( .A1(u5_mult_82_n368), .A2(u5_mult_82_n212), .ZN(
        u5_mult_82_ab_51__38_) );
  NOR2_X1 u5_mult_82_U819 ( .A1(u5_mult_82_n365), .A2(u5_mult_82_n212), .ZN(
        u5_mult_82_ab_51__39_) );
  NOR2_X1 u5_mult_82_U818 ( .A1(u5_mult_82_n441), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__3_) );
  NOR2_X1 u5_mult_82_U817 ( .A1(u5_mult_82_n363), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__40_) );
  NOR2_X1 u5_mult_82_U816 ( .A1(u5_mult_82_n361), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__41_) );
  NOR2_X1 u5_mult_82_U815 ( .A1(u5_mult_82_n360), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__42_) );
  NOR2_X1 u5_mult_82_U814 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__43_) );
  NOR2_X1 u5_mult_82_U813 ( .A1(u5_mult_82_n355), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__44_) );
  NOR2_X1 u5_mult_82_U812 ( .A1(u5_mult_82_n351), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__45_) );
  NOR2_X1 u5_mult_82_U811 ( .A1(u5_mult_82_n349), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__46_) );
  NOR2_X1 u5_mult_82_U810 ( .A1(u5_mult_82_n347), .A2(u5_mult_82_n212), .ZN(
        u5_mult_82_ab_51__47_) );
  NOR2_X1 u5_mult_82_U809 ( .A1(u5_mult_82_n345), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__48_) );
  NOR2_X1 u5_mult_82_U808 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n212), .ZN(
        u5_mult_82_ab_51__49_) );
  NOR2_X1 u5_mult_82_U807 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n212), .ZN(
        u5_mult_82_ab_51__4_) );
  NOR2_X1 u5_mult_82_U806 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__50_) );
  NOR2_X1 u5_mult_82_U805 ( .A1(u5_mult_82_n340), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__51_) );
  NOR2_X1 u5_mult_82_U804 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__52_) );
  NOR2_X1 u5_mult_82_U803 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__5_) );
  NOR2_X1 u5_mult_82_U802 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__6_) );
  NOR2_X1 u5_mult_82_U801 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__7_) );
  NOR2_X1 u5_mult_82_U800 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__8_) );
  NOR2_X1 u5_mult_82_U799 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n211), .ZN(
        u5_mult_82_ab_51__9_) );
  NOR2_X1 u5_mult_82_U798 ( .A1(u5_mult_82_n480), .A2(u5_mult_82_n447), .ZN(
        u5_mult_82_ab_52__0_) );
  NOR2_X1 u5_mult_82_U797 ( .A1(u5_mult_82_n477), .A2(u5_mult_82_n447), .ZN(
        u5_mult_82_ab_52__10_) );
  NOR2_X1 u5_mult_82_U796 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n447), .ZN(
        u5_mult_82_ab_52__11_) );
  NOR2_X1 u5_mult_82_U795 ( .A1(u5_mult_82_n424), .A2(u5_mult_82_n447), .ZN(
        u5_mult_82_ab_52__12_) );
  NOR2_X1 u5_mult_82_U794 ( .A1(u5_mult_82_n421), .A2(u5_mult_82_n447), .ZN(
        u5_mult_82_ab_52__13_) );
  NOR2_X1 u5_mult_82_U793 ( .A1(u5_mult_82_n418), .A2(u5_mult_82_n447), .ZN(
        u5_mult_82_ab_52__14_) );
  NOR2_X1 u5_mult_82_U792 ( .A1(u5_mult_82_n415), .A2(u5_mult_82_n447), .ZN(
        u5_mult_82_ab_52__15_) );
  NOR2_X1 u5_mult_82_U791 ( .A1(u5_mult_82_n412), .A2(u5_mult_82_n447), .ZN(
        u5_mult_82_ab_52__16_) );
  NOR2_X1 u5_mult_82_U790 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n447), .ZN(
        u5_mult_82_ab_52__17_) );
  NOR2_X1 u5_mult_82_U789 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n448), .ZN(
        u5_mult_82_ab_52__18_) );
  NOR2_X1 u5_mult_82_U788 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n448), .ZN(
        u5_mult_82_ab_52__19_) );
  NOR2_X1 u5_mult_82_U787 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n448), .ZN(
        u5_mult_82_ab_52__1_) );
  NOR2_X1 u5_mult_82_U786 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n448), .ZN(
        u5_mult_82_ab_52__20_) );
  NOR2_X1 u5_mult_82_U785 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n448), .ZN(
        u5_mult_82_ab_52__21_) );
  NOR2_X1 u5_mult_82_U784 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n448), .ZN(
        u5_mult_82_ab_52__22_) );
  NOR2_X1 u5_mult_82_U783 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n448), .ZN(
        u5_mult_82_ab_52__23_) );
  NOR2_X1 u5_mult_82_U782 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n448), .ZN(
        u5_mult_82_ab_52__24_) );
  NOR2_X1 u5_mult_82_U781 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n448), .ZN(
        u5_mult_82_ab_52__25_) );
  NOR2_X1 u5_mult_82_U780 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n448), .ZN(
        u5_mult_82_ab_52__26_) );
  NOR2_X1 u5_mult_82_U779 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n448), .ZN(
        u5_mult_82_ab_52__27_) );
  NOR2_X1 u5_mult_82_U778 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n449), .ZN(
        u5_mult_82_ab_52__28_) );
  NOR2_X1 u5_mult_82_U777 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n449), .ZN(
        u5_mult_82_ab_52__29_) );
  NOR2_X1 u5_mult_82_U776 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n449), .ZN(
        u5_mult_82_ab_52__2_) );
  NOR2_X1 u5_mult_82_U775 ( .A1(u5_mult_82_n384), .A2(u5_mult_82_n449), .ZN(
        u5_mult_82_ab_52__30_) );
  NOR2_X1 u5_mult_82_U774 ( .A1(u5_mult_82_n382), .A2(u5_mult_82_n448), .ZN(
        u5_mult_82_ab_52__31_) );
  NOR2_X1 u5_mult_82_U773 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n449), .ZN(
        u5_mult_82_ab_52__32_) );
  NOR2_X1 u5_mult_82_U772 ( .A1(u5_mult_82_n378), .A2(u5_mult_82_n449), .ZN(
        u5_mult_82_ab_52__33_) );
  NOR2_X1 u5_mult_82_U771 ( .A1(u5_mult_82_n376), .A2(u5_mult_82_n449), .ZN(
        u5_mult_82_ab_52__34_) );
  NOR2_X1 u5_mult_82_U770 ( .A1(u5_mult_82_n374), .A2(u5_mult_82_n449), .ZN(
        u5_mult_82_ab_52__35_) );
  NOR2_X1 u5_mult_82_U769 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n449), .ZN(
        u5_mult_82_ab_52__36_) );
  NOR2_X1 u5_mult_82_U768 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n447), .ZN(
        u5_mult_82_ab_52__37_) );
  NOR2_X1 u5_mult_82_U767 ( .A1(u5_mult_82_n368), .A2(u5_mult_82_n448), .ZN(
        u5_mult_82_ab_52__38_) );
  NOR2_X1 u5_mult_82_U766 ( .A1(u5_mult_82_n366), .A2(u5_mult_82_n448), .ZN(
        u5_mult_82_ab_52__39_) );
  NOR2_X1 u5_mult_82_U765 ( .A1(u5_mult_82_n441), .A2(u5_mult_82_n447), .ZN(
        u5_mult_82_ab_52__3_) );
  NOR2_X1 u5_mult_82_U764 ( .A1(u5_mult_82_n364), .A2(u5_mult_82_n448), .ZN(
        u5_mult_82_ab_52__40_) );
  NOR2_X1 u5_mult_82_U763 ( .A1(u5_mult_82_n362), .A2(u5_mult_82_n448), .ZN(
        u5_mult_82_ab_52__41_) );
  NOR2_X1 u5_mult_82_U762 ( .A1(u5_mult_82_n360), .A2(u5_mult_82_n448), .ZN(
        u5_mult_82_ab_52__42_) );
  NOR2_X1 u5_mult_82_U761 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n448), .ZN(
        u5_mult_82_ab_52__43_) );
  NOR2_X1 u5_mult_82_U760 ( .A1(u5_mult_82_n355), .A2(u5_mult_82_n448), .ZN(
        u5_mult_82_ab_52__44_) );
  NOR2_X1 u5_mult_82_U759 ( .A1(u5_mult_82_n352), .A2(u5_mult_82_n448), .ZN(
        u5_mult_82_ab_52__45_) );
  NOR2_X1 u5_mult_82_U758 ( .A1(u5_mult_82_n350), .A2(u5_mult_82_n448), .ZN(
        u5_mult_82_ab_52__46_) );
  NOR2_X1 u5_mult_82_U757 ( .A1(u5_mult_82_n348), .A2(u5_mult_82_n448), .ZN(
        u5_mult_82_ab_52__47_) );
  NOR2_X1 u5_mult_82_U756 ( .A1(u5_mult_82_n346), .A2(u5_mult_82_n447), .ZN(
        u5_mult_82_ab_52__48_) );
  NOR2_X1 u5_mult_82_U755 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n447), .ZN(
        u5_mult_82_ab_52__49_) );
  NOR2_X1 u5_mult_82_U754 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n447), .ZN(
        u5_mult_82_ab_52__4_) );
  NOR2_X1 u5_mult_82_U753 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n447), .ZN(
        u5_mult_82_ab_52__50_) );
  NOR2_X1 u5_mult_82_U752 ( .A1(u5_mult_82_n340), .A2(u5_mult_82_n447), .ZN(
        u5_mult_82_ab_52__51_) );
  NOR2_X1 u5_mult_82_U751 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n447), .ZN(
        u5_mult_82_ab_52__52_) );
  NOR2_X1 u5_mult_82_U750 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n447), .ZN(
        u5_mult_82_ab_52__5_) );
  NOR2_X1 u5_mult_82_U749 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n447), .ZN(
        u5_mult_82_ab_52__6_) );
  NOR2_X1 u5_mult_82_U748 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n447), .ZN(
        u5_mult_82_ab_52__7_) );
  NOR2_X1 u5_mult_82_U747 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n447), .ZN(
        u5_mult_82_ab_52__8_) );
  NOR2_X1 u5_mult_82_U746 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n447), .ZN(
        u5_mult_82_ab_52__9_) );
  NOR2_X1 u5_mult_82_U745 ( .A1(u5_mult_82_n480), .A2(u5_mult_82_n319), .ZN(
        u5_mult_82_ab_5__0_) );
  NOR2_X1 u5_mult_82_U744 ( .A1(u5_mult_82_n477), .A2(u5_mult_82_n319), .ZN(
        u5_mult_82_ab_5__10_) );
  NOR2_X1 u5_mult_82_U743 ( .A1(u5_mult_82_n426), .A2(u5_mult_82_n319), .ZN(
        u5_mult_82_ab_5__11_) );
  NOR2_X1 u5_mult_82_U742 ( .A1(u5_mult_82_n424), .A2(u5_mult_82_n319), .ZN(
        u5_mult_82_ab_5__12_) );
  NOR2_X1 u5_mult_82_U741 ( .A1(u5_mult_82_n421), .A2(u5_mult_82_n319), .ZN(
        u5_mult_82_ab_5__13_) );
  NOR2_X1 u5_mult_82_U740 ( .A1(u5_mult_82_n418), .A2(u5_mult_82_n319), .ZN(
        u5_mult_82_ab_5__14_) );
  NOR2_X1 u5_mult_82_U739 ( .A1(u5_mult_82_n415), .A2(u5_mult_82_n319), .ZN(
        u5_mult_82_ab_5__15_) );
  NOR2_X1 u5_mult_82_U738 ( .A1(u5_mult_82_n412), .A2(u5_mult_82_n319), .ZN(
        u5_mult_82_ab_5__16_) );
  NOR2_X1 u5_mult_82_U737 ( .A1(u5_mult_82_n409), .A2(u5_mult_82_n319), .ZN(
        u5_mult_82_ab_5__17_) );
  NOR2_X1 u5_mult_82_U736 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n319), .ZN(
        u5_mult_82_ab_5__18_) );
  NOR2_X1 u5_mult_82_U735 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n319), .ZN(
        u5_mult_82_ab_5__19_) );
  NOR2_X1 u5_mult_82_U734 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n320), .ZN(
        u5_mult_82_ab_5__1_) );
  NOR2_X1 u5_mult_82_U733 ( .A1(u5_mult_82_n475), .A2(u5_mult_82_n320), .ZN(
        u5_mult_82_ab_5__20_) );
  NOR2_X1 u5_mult_82_U732 ( .A1(u5_mult_82_n402), .A2(u5_mult_82_n320), .ZN(
        u5_mult_82_ab_5__21_) );
  NOR2_X1 u5_mult_82_U731 ( .A1(u5_mult_82_n400), .A2(u5_mult_82_n320), .ZN(
        u5_mult_82_ab_5__22_) );
  NOR2_X1 u5_mult_82_U730 ( .A1(u5_mult_82_n398), .A2(u5_mult_82_n320), .ZN(
        u5_mult_82_ab_5__23_) );
  NOR2_X1 u5_mult_82_U729 ( .A1(u5_mult_82_n396), .A2(u5_mult_82_n320), .ZN(
        u5_mult_82_ab_5__24_) );
  NOR2_X1 u5_mult_82_U728 ( .A1(u5_mult_82_n394), .A2(u5_mult_82_n320), .ZN(
        u5_mult_82_ab_5__25_) );
  NOR2_X1 u5_mult_82_U727 ( .A1(u5_mult_82_n392), .A2(u5_mult_82_n320), .ZN(
        u5_mult_82_ab_5__26_) );
  NOR2_X1 u5_mult_82_U726 ( .A1(u5_mult_82_n390), .A2(u5_mult_82_n320), .ZN(
        u5_mult_82_ab_5__27_) );
  NOR2_X1 u5_mult_82_U725 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n320), .ZN(
        u5_mult_82_ab_5__28_) );
  NOR2_X1 u5_mult_82_U724 ( .A1(u5_mult_82_n386), .A2(u5_mult_82_n320), .ZN(
        u5_mult_82_ab_5__29_) );
  NOR2_X1 u5_mult_82_U723 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n321), .ZN(
        u5_mult_82_ab_5__2_) );
  NOR2_X1 u5_mult_82_U722 ( .A1(u5_mult_82_n384), .A2(u5_mult_82_n321), .ZN(
        u5_mult_82_ab_5__30_) );
  NOR2_X1 u5_mult_82_U721 ( .A1(u5_mult_82_n382), .A2(u5_mult_82_n321), .ZN(
        u5_mult_82_ab_5__31_) );
  NOR2_X1 u5_mult_82_U720 ( .A1(u5_mult_82_n380), .A2(u5_mult_82_n321), .ZN(
        u5_mult_82_ab_5__32_) );
  NOR2_X1 u5_mult_82_U719 ( .A1(u5_mult_82_n378), .A2(u5_mult_82_n321), .ZN(
        u5_mult_82_ab_5__33_) );
  NOR2_X1 u5_mult_82_U718 ( .A1(u5_mult_82_n376), .A2(u5_mult_82_n321), .ZN(
        u5_mult_82_ab_5__34_) );
  NOR2_X1 u5_mult_82_U717 ( .A1(u5_mult_82_n374), .A2(u5_mult_82_n321), .ZN(
        u5_mult_82_ab_5__35_) );
  NOR2_X1 u5_mult_82_U716 ( .A1(u5_mult_82_n474), .A2(u5_mult_82_n321), .ZN(
        u5_mult_82_ab_5__36_) );
  NOR2_X1 u5_mult_82_U715 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n321), .ZN(
        u5_mult_82_ab_5__37_) );
  NOR2_X1 u5_mult_82_U714 ( .A1(u5_mult_82_n368), .A2(u5_mult_82_n321), .ZN(
        u5_mult_82_ab_5__38_) );
  NOR2_X1 u5_mult_82_U713 ( .A1(u5_mult_82_n366), .A2(u5_mult_82_n321), .ZN(
        u5_mult_82_ab_5__39_) );
  NOR2_X1 u5_mult_82_U712 ( .A1(u5_mult_82_n441), .A2(u5_mult_82_n319), .ZN(
        u5_mult_82_ab_5__3_) );
  NOR2_X1 u5_mult_82_U711 ( .A1(u5_mult_82_n364), .A2(u5_mult_82_n319), .ZN(
        u5_mult_82_ab_5__40_) );
  NOR2_X1 u5_mult_82_U710 ( .A1(u5_mult_82_n362), .A2(u5_mult_82_n320), .ZN(
        u5_mult_82_ab_5__41_) );
  NOR2_X1 u5_mult_82_U709 ( .A1(u5_mult_82_n360), .A2(u5_mult_82_n321), .ZN(
        u5_mult_82_ab_5__42_) );
  NOR2_X1 u5_mult_82_U708 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n320), .ZN(
        u5_mult_82_ab_5__43_) );
  NOR2_X1 u5_mult_82_U707 ( .A1(u5_mult_82_n355), .A2(u5_mult_82_n321), .ZN(
        u5_mult_82_ab_5__44_) );
  NOR2_X1 u5_mult_82_U706 ( .A1(u5_mult_82_n352), .A2(u5_mult_82_n320), .ZN(
        u5_mult_82_ab_5__45_) );
  NOR2_X1 u5_mult_82_U705 ( .A1(u5_mult_82_n350), .A2(u5_mult_82_n319), .ZN(
        u5_mult_82_ab_5__46_) );
  NOR2_X1 u5_mult_82_U704 ( .A1(u5_mult_82_n348), .A2(u5_mult_82_n319), .ZN(
        u5_mult_82_ab_5__47_) );
  NOR2_X1 u5_mult_82_U703 ( .A1(u5_mult_82_n346), .A2(u5_mult_82_n322), .ZN(
        u5_mult_82_ab_5__48_) );
  NOR2_X1 u5_mult_82_U702 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n322), .ZN(
        u5_mult_82_ab_5__49_) );
  NOR2_X1 u5_mult_82_U701 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n319), .ZN(
        u5_mult_82_ab_5__4_) );
  NOR2_X1 u5_mult_82_U700 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n322), .ZN(
        u5_mult_82_ab_5__50_) );
  NOR2_X1 u5_mult_82_U699 ( .A1(u5_mult_82_n340), .A2(u5_mult_82_n321), .ZN(
        u5_mult_82_ab_5__51_) );
  NOR2_X1 u5_mult_82_U698 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n320), .ZN(
        u5_mult_82_ab_5__52_) );
  NOR2_X1 u5_mult_82_U697 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n319), .ZN(
        u5_mult_82_ab_5__5_) );
  NOR2_X1 u5_mult_82_U696 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n319), .ZN(
        u5_mult_82_ab_5__6_) );
  NOR2_X1 u5_mult_82_U695 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n319), .ZN(
        u5_mult_82_ab_5__7_) );
  NOR2_X1 u5_mult_82_U694 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n319), .ZN(
        u5_mult_82_ab_5__8_) );
  NOR2_X1 u5_mult_82_U693 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n319), .ZN(
        u5_mult_82_ab_5__9_) );
  NOR2_X1 u5_mult_82_U692 ( .A1(u5_mult_82_n480), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__0_) );
  NOR2_X1 u5_mult_82_U691 ( .A1(u5_mult_82_n477), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__10_) );
  NOR2_X1 u5_mult_82_U690 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__11_) );
  NOR2_X1 u5_mult_82_U689 ( .A1(u5_mult_82_n424), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__12_) );
  NOR2_X1 u5_mult_82_U688 ( .A1(u5_mult_82_n421), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__13_) );
  NOR2_X1 u5_mult_82_U687 ( .A1(u5_mult_82_n418), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__14_) );
  NOR2_X1 u5_mult_82_U686 ( .A1(u5_mult_82_n415), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__15_) );
  NOR2_X1 u5_mult_82_U685 ( .A1(u5_mult_82_n412), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__16_) );
  NOR2_X1 u5_mult_82_U684 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__17_) );
  NOR2_X1 u5_mult_82_U683 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__18_) );
  NOR2_X1 u5_mult_82_U682 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__19_) );
  NOR2_X1 u5_mult_82_U681 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__1_) );
  NOR2_X1 u5_mult_82_U680 ( .A1(u5_mult_82_n475), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__20_) );
  NOR2_X1 u5_mult_82_U679 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__21_) );
  NOR2_X1 u5_mult_82_U678 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__22_) );
  NOR2_X1 u5_mult_82_U677 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__23_) );
  NOR2_X1 u5_mult_82_U676 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__24_) );
  NOR2_X1 u5_mult_82_U675 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__25_) );
  NOR2_X1 u5_mult_82_U674 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__26_) );
  NOR2_X1 u5_mult_82_U673 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__27_) );
  NOR2_X1 u5_mult_82_U672 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__28_) );
  NOR2_X1 u5_mult_82_U671 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__29_) );
  NOR2_X1 u5_mult_82_U670 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n317), .ZN(
        u5_mult_82_ab_6__2_) );
  NOR2_X1 u5_mult_82_U669 ( .A1(u5_mult_82_n384), .A2(u5_mult_82_n317), .ZN(
        u5_mult_82_ab_6__30_) );
  NOR2_X1 u5_mult_82_U668 ( .A1(u5_mult_82_n382), .A2(u5_mult_82_n317), .ZN(
        u5_mult_82_ab_6__31_) );
  NOR2_X1 u5_mult_82_U667 ( .A1(u5_mult_82_n380), .A2(u5_mult_82_n317), .ZN(
        u5_mult_82_ab_6__32_) );
  NOR2_X1 u5_mult_82_U666 ( .A1(u5_mult_82_n378), .A2(u5_mult_82_n317), .ZN(
        u5_mult_82_ab_6__33_) );
  NOR2_X1 u5_mult_82_U665 ( .A1(u5_mult_82_n376), .A2(u5_mult_82_n317), .ZN(
        u5_mult_82_ab_6__34_) );
  NOR2_X1 u5_mult_82_U664 ( .A1(u5_mult_82_n374), .A2(u5_mult_82_n317), .ZN(
        u5_mult_82_ab_6__35_) );
  NOR2_X1 u5_mult_82_U663 ( .A1(u5_mult_82_n474), .A2(u5_mult_82_n317), .ZN(
        u5_mult_82_ab_6__36_) );
  NOR2_X1 u5_mult_82_U662 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n317), .ZN(
        u5_mult_82_ab_6__37_) );
  NOR2_X1 u5_mult_82_U661 ( .A1(u5_mult_82_n368), .A2(u5_mult_82_n317), .ZN(
        u5_mult_82_ab_6__38_) );
  NOR2_X1 u5_mult_82_U660 ( .A1(u5_mult_82_n366), .A2(u5_mult_82_n317), .ZN(
        u5_mult_82_ab_6__39_) );
  NOR2_X1 u5_mult_82_U659 ( .A1(u5_mult_82_n441), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__3_) );
  NOR2_X1 u5_mult_82_U658 ( .A1(u5_mult_82_n364), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__40_) );
  NOR2_X1 u5_mult_82_U657 ( .A1(u5_mult_82_n362), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__41_) );
  NOR2_X1 u5_mult_82_U656 ( .A1(u5_mult_82_n360), .A2(u5_mult_82_n318), .ZN(
        u5_mult_82_ab_6__42_) );
  NOR2_X1 u5_mult_82_U655 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n318), .ZN(
        u5_mult_82_ab_6__43_) );
  NOR2_X1 u5_mult_82_U654 ( .A1(u5_mult_82_n355), .A2(u5_mult_82_n318), .ZN(
        u5_mult_82_ab_6__44_) );
  NOR2_X1 u5_mult_82_U653 ( .A1(u5_mult_82_n352), .A2(u5_mult_82_n317), .ZN(
        u5_mult_82_ab_6__45_) );
  NOR2_X1 u5_mult_82_U652 ( .A1(u5_mult_82_n350), .A2(u5_mult_82_n318), .ZN(
        u5_mult_82_ab_6__46_) );
  NOR2_X1 u5_mult_82_U651 ( .A1(u5_mult_82_n348), .A2(u5_mult_82_n318), .ZN(
        u5_mult_82_ab_6__47_) );
  NOR2_X1 u5_mult_82_U650 ( .A1(u5_mult_82_n346), .A2(u5_mult_82_n318), .ZN(
        u5_mult_82_ab_6__48_) );
  NOR2_X1 u5_mult_82_U649 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n318), .ZN(
        u5_mult_82_ab_6__49_) );
  NOR2_X1 u5_mult_82_U648 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__4_) );
  NOR2_X1 u5_mult_82_U647 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n317), .ZN(
        u5_mult_82_ab_6__50_) );
  NOR2_X1 u5_mult_82_U646 ( .A1(u5_mult_82_n340), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__51_) );
  NOR2_X1 u5_mult_82_U645 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__52_) );
  NOR2_X1 u5_mult_82_U644 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__5_) );
  NOR2_X1 u5_mult_82_U643 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__6_) );
  NOR2_X1 u5_mult_82_U642 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__7_) );
  NOR2_X1 u5_mult_82_U641 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__8_) );
  NOR2_X1 u5_mult_82_U640 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n316), .ZN(
        u5_mult_82_ab_6__9_) );
  NOR2_X1 u5_mult_82_U639 ( .A1(u5_mult_82_n480), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__0_) );
  NOR2_X1 u5_mult_82_U638 ( .A1(u5_mult_82_n477), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__10_) );
  NOR2_X1 u5_mult_82_U637 ( .A1(u5_mult_82_n426), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__11_) );
  NOR2_X1 u5_mult_82_U636 ( .A1(u5_mult_82_n424), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__12_) );
  NOR2_X1 u5_mult_82_U635 ( .A1(u5_mult_82_n421), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__13_) );
  NOR2_X1 u5_mult_82_U634 ( .A1(u5_mult_82_n418), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__14_) );
  NOR2_X1 u5_mult_82_U633 ( .A1(u5_mult_82_n415), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__15_) );
  NOR2_X1 u5_mult_82_U632 ( .A1(u5_mult_82_n412), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__16_) );
  NOR2_X1 u5_mult_82_U631 ( .A1(u5_mult_82_n409), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__17_) );
  NOR2_X1 u5_mult_82_U630 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__18_) );
  NOR2_X1 u5_mult_82_U629 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__19_) );
  NOR2_X1 u5_mult_82_U628 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n315), .ZN(
        u5_mult_82_ab_7__1_) );
  NOR2_X1 u5_mult_82_U627 ( .A1(u5_mult_82_n403), .A2(u5_mult_82_n315), .ZN(
        u5_mult_82_ab_7__20_) );
  NOR2_X1 u5_mult_82_U626 ( .A1(u5_mult_82_n402), .A2(u5_mult_82_n315), .ZN(
        u5_mult_82_ab_7__21_) );
  NOR2_X1 u5_mult_82_U625 ( .A1(u5_mult_82_n400), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__22_) );
  NOR2_X1 u5_mult_82_U624 ( .A1(u5_mult_82_n398), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__23_) );
  NOR2_X1 u5_mult_82_U623 ( .A1(u5_mult_82_n396), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__24_) );
  NOR2_X1 u5_mult_82_U622 ( .A1(u5_mult_82_n394), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__25_) );
  NOR2_X1 u5_mult_82_U621 ( .A1(u5_mult_82_n392), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__26_) );
  NOR2_X1 u5_mult_82_U620 ( .A1(u5_mult_82_n390), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__27_) );
  NOR2_X1 u5_mult_82_U619 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__28_) );
  NOR2_X1 u5_mult_82_U618 ( .A1(u5_mult_82_n386), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__29_) );
  NOR2_X1 u5_mult_82_U617 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n315), .ZN(
        u5_mult_82_ab_7__2_) );
  NOR2_X1 u5_mult_82_U616 ( .A1(u5_mult_82_n384), .A2(u5_mult_82_n315), .ZN(
        u5_mult_82_ab_7__30_) );
  NOR2_X1 u5_mult_82_U615 ( .A1(u5_mult_82_n382), .A2(u5_mult_82_n315), .ZN(
        u5_mult_82_ab_7__31_) );
  NOR2_X1 u5_mult_82_U614 ( .A1(u5_mult_82_n380), .A2(u5_mult_82_n315), .ZN(
        u5_mult_82_ab_7__32_) );
  NOR2_X1 u5_mult_82_U613 ( .A1(u5_mult_82_n378), .A2(u5_mult_82_n315), .ZN(
        u5_mult_82_ab_7__33_) );
  NOR2_X1 u5_mult_82_U612 ( .A1(u5_mult_82_n376), .A2(u5_mult_82_n315), .ZN(
        u5_mult_82_ab_7__34_) );
  NOR2_X1 u5_mult_82_U611 ( .A1(u5_mult_82_n374), .A2(u5_mult_82_n315), .ZN(
        u5_mult_82_ab_7__35_) );
  NOR2_X1 u5_mult_82_U610 ( .A1(u5_mult_82_n474), .A2(u5_mult_82_n315), .ZN(
        u5_mult_82_ab_7__36_) );
  NOR2_X1 u5_mult_82_U609 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n315), .ZN(
        u5_mult_82_ab_7__37_) );
  NOR2_X1 u5_mult_82_U608 ( .A1(u5_mult_82_n368), .A2(u5_mult_82_n315), .ZN(
        u5_mult_82_ab_7__38_) );
  NOR2_X1 u5_mult_82_U607 ( .A1(u5_mult_82_n366), .A2(u5_mult_82_n315), .ZN(
        u5_mult_82_ab_7__39_) );
  NOR2_X1 u5_mult_82_U606 ( .A1(u5_mult_82_n441), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__3_) );
  NOR2_X1 u5_mult_82_U605 ( .A1(u5_mult_82_n364), .A2(u5_mult_82_n473), .ZN(
        u5_mult_82_ab_7__40_) );
  NOR2_X1 u5_mult_82_U604 ( .A1(u5_mult_82_n362), .A2(u5_mult_82_n473), .ZN(
        u5_mult_82_ab_7__41_) );
  NOR2_X1 u5_mult_82_U603 ( .A1(u5_mult_82_n360), .A2(u5_mult_82_n315), .ZN(
        u5_mult_82_ab_7__42_) );
  NOR2_X1 u5_mult_82_U602 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n315), .ZN(
        u5_mult_82_ab_7__43_) );
  NOR2_X1 u5_mult_82_U601 ( .A1(u5_mult_82_n355), .A2(u5_mult_82_n473), .ZN(
        u5_mult_82_ab_7__44_) );
  NOR2_X1 u5_mult_82_U600 ( .A1(u5_mult_82_n352), .A2(u5_mult_82_n473), .ZN(
        u5_mult_82_ab_7__45_) );
  NOR2_X1 u5_mult_82_U599 ( .A1(u5_mult_82_n350), .A2(u5_mult_82_n473), .ZN(
        u5_mult_82_ab_7__46_) );
  NOR2_X1 u5_mult_82_U598 ( .A1(u5_mult_82_n348), .A2(u5_mult_82_n473), .ZN(
        u5_mult_82_ab_7__47_) );
  NOR2_X1 u5_mult_82_U597 ( .A1(u5_mult_82_n346), .A2(u5_mult_82_n473), .ZN(
        u5_mult_82_ab_7__48_) );
  NOR2_X1 u5_mult_82_U596 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n315), .ZN(
        u5_mult_82_ab_7__49_) );
  NOR2_X1 u5_mult_82_U595 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__4_) );
  NOR2_X1 u5_mult_82_U594 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__50_) );
  NOR2_X1 u5_mult_82_U593 ( .A1(u5_mult_82_n340), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__51_) );
  NOR2_X1 u5_mult_82_U592 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__52_) );
  NOR2_X1 u5_mult_82_U591 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__5_) );
  NOR2_X1 u5_mult_82_U590 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__6_) );
  NOR2_X1 u5_mult_82_U589 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__7_) );
  NOR2_X1 u5_mult_82_U588 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__8_) );
  NOR2_X1 u5_mult_82_U587 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n314), .ZN(
        u5_mult_82_ab_7__9_) );
  NOR2_X1 u5_mult_82_U586 ( .A1(u5_mult_82_n480), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__0_) );
  NOR2_X1 u5_mult_82_U585 ( .A1(u5_mult_82_n427), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__10_) );
  NOR2_X1 u5_mult_82_U584 ( .A1(u5_mult_82_n425), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__11_) );
  NOR2_X1 u5_mult_82_U583 ( .A1(u5_mult_82_n424), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__12_) );
  NOR2_X1 u5_mult_82_U582 ( .A1(u5_mult_82_n421), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__13_) );
  NOR2_X1 u5_mult_82_U581 ( .A1(u5_mult_82_n418), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__14_) );
  NOR2_X1 u5_mult_82_U580 ( .A1(u5_mult_82_n415), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__15_) );
  NOR2_X1 u5_mult_82_U579 ( .A1(u5_mult_82_n412), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__16_) );
  NOR2_X1 u5_mult_82_U578 ( .A1(u5_mult_82_n408), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__17_) );
  NOR2_X1 u5_mult_82_U577 ( .A1(u5_mult_82_n407), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__18_) );
  NOR2_X1 u5_mult_82_U576 ( .A1(u5_mult_82_n405), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__19_) );
  NOR2_X1 u5_mult_82_U575 ( .A1(u5_mult_82_n444), .A2(u5_mult_82_n313), .ZN(
        u5_mult_82_ab_8__1_) );
  NOR2_X1 u5_mult_82_U574 ( .A1(u5_mult_82_n475), .A2(u5_mult_82_n313), .ZN(
        u5_mult_82_ab_8__20_) );
  NOR2_X1 u5_mult_82_U573 ( .A1(u5_mult_82_n401), .A2(u5_mult_82_n313), .ZN(
        u5_mult_82_ab_8__21_) );
  NOR2_X1 u5_mult_82_U572 ( .A1(u5_mult_82_n399), .A2(u5_mult_82_n313), .ZN(
        u5_mult_82_ab_8__22_) );
  NOR2_X1 u5_mult_82_U571 ( .A1(u5_mult_82_n397), .A2(u5_mult_82_n313), .ZN(
        u5_mult_82_ab_8__23_) );
  NOR2_X1 u5_mult_82_U570 ( .A1(u5_mult_82_n395), .A2(u5_mult_82_n313), .ZN(
        u5_mult_82_ab_8__24_) );
  NOR2_X1 u5_mult_82_U569 ( .A1(u5_mult_82_n393), .A2(u5_mult_82_n313), .ZN(
        u5_mult_82_ab_8__25_) );
  NOR2_X1 u5_mult_82_U568 ( .A1(u5_mult_82_n391), .A2(u5_mult_82_n313), .ZN(
        u5_mult_82_ab_8__26_) );
  NOR2_X1 u5_mult_82_U567 ( .A1(u5_mult_82_n389), .A2(u5_mult_82_n313), .ZN(
        u5_mult_82_ab_8__27_) );
  NOR2_X1 u5_mult_82_U566 ( .A1(u5_mult_82_n388), .A2(u5_mult_82_n313), .ZN(
        u5_mult_82_ab_8__28_) );
  NOR2_X1 u5_mult_82_U565 ( .A1(u5_mult_82_n385), .A2(u5_mult_82_n313), .ZN(
        u5_mult_82_ab_8__29_) );
  NOR2_X1 u5_mult_82_U564 ( .A1(u5_mult_82_n479), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__2_) );
  NOR2_X1 u5_mult_82_U563 ( .A1(u5_mult_82_n384), .A2(u5_mult_82_n313), .ZN(
        u5_mult_82_ab_8__30_) );
  NOR2_X1 u5_mult_82_U562 ( .A1(u5_mult_82_n382), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__31_) );
  NOR2_X1 u5_mult_82_U561 ( .A1(u5_mult_82_n379), .A2(u5_mult_82_n313), .ZN(
        u5_mult_82_ab_8__32_) );
  NOR2_X1 u5_mult_82_U560 ( .A1(u5_mult_82_n378), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__33_) );
  NOR2_X1 u5_mult_82_U559 ( .A1(u5_mult_82_n376), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__34_) );
  NOR2_X1 u5_mult_82_U558 ( .A1(u5_mult_82_n374), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__35_) );
  NOR2_X1 u5_mult_82_U557 ( .A1(u5_mult_82_n372), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__36_) );
  NOR2_X1 u5_mult_82_U556 ( .A1(u5_mult_82_n371), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__37_) );
  NOR2_X1 u5_mult_82_U555 ( .A1(u5_mult_82_n368), .A2(u5_mult_82_n313), .ZN(
        u5_mult_82_ab_8__38_) );
  NOR2_X1 u5_mult_82_U554 ( .A1(u5_mult_82_n366), .A2(u5_mult_82_n313), .ZN(
        u5_mult_82_ab_8__39_) );
  NOR2_X1 u5_mult_82_U553 ( .A1(u5_mult_82_n441), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__3_) );
  NOR2_X1 u5_mult_82_U552 ( .A1(u5_mult_82_n364), .A2(u5_mult_82_n472), .ZN(
        u5_mult_82_ab_8__40_) );
  NOR2_X1 u5_mult_82_U551 ( .A1(u5_mult_82_n362), .A2(u5_mult_82_n313), .ZN(
        u5_mult_82_ab_8__41_) );
  NOR2_X1 u5_mult_82_U550 ( .A1(u5_mult_82_n360), .A2(u5_mult_82_n472), .ZN(
        u5_mult_82_ab_8__42_) );
  NOR2_X1 u5_mult_82_U549 ( .A1(u5_mult_82_n357), .A2(u5_mult_82_n472), .ZN(
        u5_mult_82_ab_8__43_) );
  NOR2_X1 u5_mult_82_U548 ( .A1(u5_mult_82_n355), .A2(u5_mult_82_n472), .ZN(
        u5_mult_82_ab_8__44_) );
  NOR2_X1 u5_mult_82_U547 ( .A1(u5_mult_82_n352), .A2(u5_mult_82_n472), .ZN(
        u5_mult_82_ab_8__45_) );
  NOR2_X1 u5_mult_82_U546 ( .A1(u5_mult_82_n350), .A2(u5_mult_82_n472), .ZN(
        u5_mult_82_ab_8__46_) );
  NOR2_X1 u5_mult_82_U545 ( .A1(u5_mult_82_n348), .A2(u5_mult_82_n472), .ZN(
        u5_mult_82_ab_8__47_) );
  NOR2_X1 u5_mult_82_U544 ( .A1(u5_mult_82_n346), .A2(u5_mult_82_n472), .ZN(
        u5_mult_82_ab_8__48_) );
  NOR2_X1 u5_mult_82_U543 ( .A1(u5_mult_82_n344), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__49_) );
  NOR2_X1 u5_mult_82_U542 ( .A1(u5_mult_82_n439), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__4_) );
  NOR2_X1 u5_mult_82_U541 ( .A1(u5_mult_82_n341), .A2(u5_mult_82_n313), .ZN(
        u5_mult_82_ab_8__50_) );
  NOR2_X1 u5_mult_82_U540 ( .A1(u5_mult_82_n340), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__51_) );
  NOR2_X1 u5_mult_82_U539 ( .A1(u5_mult_82_n337), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__52_) );
  NOR2_X1 u5_mult_82_U538 ( .A1(u5_mult_82_n437), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__5_) );
  NOR2_X1 u5_mult_82_U537 ( .A1(u5_mult_82_n435), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__6_) );
  NOR2_X1 u5_mult_82_U536 ( .A1(u5_mult_82_n433), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__7_) );
  NOR2_X1 u5_mult_82_U535 ( .A1(u5_mult_82_n431), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__8_) );
  NOR2_X1 u5_mult_82_U534 ( .A1(u5_mult_82_n429), .A2(u5_mult_82_n312), .ZN(
        u5_mult_82_ab_8__9_) );
  NOR2_X1 u5_mult_82_U533 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n446), .ZN(
        u5_mult_82_ab_9__0_) );
  NOR2_X1 u5_mult_82_U532 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n477), .ZN(
        u5_mult_82_ab_9__10_) );
  NOR2_X1 u5_mult_82_U531 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n426), .ZN(
        u5_mult_82_ab_9__11_) );
  NOR2_X1 u5_mult_82_U530 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n424), .ZN(
        u5_mult_82_ab_9__12_) );
  NOR2_X1 u5_mult_82_U529 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n421), .ZN(
        u5_mult_82_ab_9__13_) );
  NOR2_X1 u5_mult_82_U528 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n418), .ZN(
        u5_mult_82_ab_9__14_) );
  NOR2_X1 u5_mult_82_U527 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n415), .ZN(
        u5_mult_82_ab_9__15_) );
  NOR2_X1 u5_mult_82_U526 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n412), .ZN(
        u5_mult_82_ab_9__16_) );
  NOR2_X1 u5_mult_82_U525 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n409), .ZN(
        u5_mult_82_ab_9__17_) );
  NOR2_X1 u5_mult_82_U524 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n407), .ZN(
        u5_mult_82_ab_9__18_) );
  NOR2_X1 u5_mult_82_U523 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n405), .ZN(
        u5_mult_82_ab_9__19_) );
  NOR2_X1 u5_mult_82_U522 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n444), .ZN(
        u5_mult_82_ab_9__1_) );
  NOR2_X1 u5_mult_82_U521 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n475), .ZN(
        u5_mult_82_ab_9__20_) );
  NOR2_X1 u5_mult_82_U520 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n402), .ZN(
        u5_mult_82_ab_9__21_) );
  NOR2_X1 u5_mult_82_U519 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n400), .ZN(
        u5_mult_82_ab_9__22_) );
  NOR2_X1 u5_mult_82_U518 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n398), .ZN(
        u5_mult_82_ab_9__23_) );
  NOR2_X1 u5_mult_82_U517 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n396), .ZN(
        u5_mult_82_ab_9__24_) );
  NOR2_X1 u5_mult_82_U516 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n394), .ZN(
        u5_mult_82_ab_9__25_) );
  NOR2_X1 u5_mult_82_U515 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n392), .ZN(
        u5_mult_82_ab_9__26_) );
  NOR2_X1 u5_mult_82_U514 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n390), .ZN(
        u5_mult_82_ab_9__27_) );
  NOR2_X1 u5_mult_82_U513 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n388), .ZN(
        u5_mult_82_ab_9__28_) );
  NOR2_X1 u5_mult_82_U512 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n386), .ZN(
        u5_mult_82_ab_9__29_) );
  NOR2_X1 u5_mult_82_U511 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n479), .ZN(
        u5_mult_82_ab_9__2_) );
  NOR2_X1 u5_mult_82_U510 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n383), .ZN(
        u5_mult_82_ab_9__30_) );
  NOR2_X1 u5_mult_82_U509 ( .A1(u5_mult_82_n311), .A2(u5_mult_82_n381), .ZN(
        u5_mult_82_ab_9__31_) );
  NOR2_X1 u5_mult_82_U508 ( .A1(u5_mult_82_n311), .A2(u5_mult_82_n380), .ZN(
        u5_mult_82_ab_9__32_) );
  NOR2_X1 u5_mult_82_U507 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n377), .ZN(
        u5_mult_82_ab_9__33_) );
  NOR2_X1 u5_mult_82_U506 ( .A1(u5_mult_82_n311), .A2(u5_mult_82_n375), .ZN(
        u5_mult_82_ab_9__34_) );
  NOR2_X1 u5_mult_82_U505 ( .A1(u5_mult_82_n311), .A2(u5_mult_82_n373), .ZN(
        u5_mult_82_ab_9__35_) );
  NOR2_X1 u5_mult_82_U504 ( .A1(u5_mult_82_n311), .A2(u5_mult_82_n474), .ZN(
        u5_mult_82_ab_9__36_) );
  NOR2_X1 u5_mult_82_U503 ( .A1(u5_mult_82_n311), .A2(u5_mult_82_n371), .ZN(
        u5_mult_82_ab_9__37_) );
  NOR2_X1 u5_mult_82_U502 ( .A1(u5_mult_82_n311), .A2(u5_mult_82_n368), .ZN(
        u5_mult_82_ab_9__38_) );
  NOR2_X1 u5_mult_82_U501 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n365), .ZN(
        u5_mult_82_ab_9__39_) );
  NOR2_X1 u5_mult_82_U500 ( .A1(u5_mult_82_n311), .A2(u5_mult_82_n441), .ZN(
        u5_mult_82_ab_9__3_) );
  NOR2_X1 u5_mult_82_U499 ( .A1(u5_mult_82_n311), .A2(u5_mult_82_n363), .ZN(
        u5_mult_82_ab_9__40_) );
  NOR2_X1 u5_mult_82_U498 ( .A1(u5_mult_82_n311), .A2(u5_mult_82_n361), .ZN(
        u5_mult_82_ab_9__41_) );
  NOR2_X1 u5_mult_82_U497 ( .A1(u5_mult_82_n311), .A2(u5_mult_82_n360), .ZN(
        u5_mult_82_ab_9__42_) );
  NOR2_X1 u5_mult_82_U496 ( .A1(u5_mult_82_n311), .A2(u5_mult_82_n357), .ZN(
        u5_mult_82_ab_9__43_) );
  NOR2_X1 u5_mult_82_U495 ( .A1(u5_mult_82_n311), .A2(u5_mult_82_n355), .ZN(
        u5_mult_82_ab_9__44_) );
  NOR2_X1 u5_mult_82_U494 ( .A1(u5_mult_82_n311), .A2(u5_mult_82_n351), .ZN(
        u5_mult_82_ab_9__45_) );
  NOR2_X1 u5_mult_82_U493 ( .A1(u5_mult_82_n311), .A2(u5_mult_82_n349), .ZN(
        u5_mult_82_ab_9__46_) );
  NOR2_X1 u5_mult_82_U492 ( .A1(u5_mult_82_n311), .A2(u5_mult_82_n347), .ZN(
        u5_mult_82_ab_9__47_) );
  NOR2_X1 u5_mult_82_U491 ( .A1(u5_mult_82_n311), .A2(u5_mult_82_n345), .ZN(
        u5_mult_82_ab_9__48_) );
  NOR2_X1 u5_mult_82_U490 ( .A1(u5_mult_82_n311), .A2(u5_mult_82_n344), .ZN(
        u5_mult_82_ab_9__49_) );
  NOR2_X1 u5_mult_82_U489 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n439), .ZN(
        u5_mult_82_ab_9__4_) );
  NOR2_X1 u5_mult_82_U488 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n341), .ZN(
        u5_mult_82_ab_9__50_) );
  NOR2_X1 u5_mult_82_U487 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n340), .ZN(
        u5_mult_82_ab_9__51_) );
  NOR2_X1 u5_mult_82_U486 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n337), .ZN(
        u5_mult_82_ab_9__52_) );
  NOR2_X1 u5_mult_82_U485 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n437), .ZN(
        u5_mult_82_ab_9__5_) );
  NOR2_X1 u5_mult_82_U484 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n435), .ZN(
        u5_mult_82_ab_9__6_) );
  NOR2_X1 u5_mult_82_U483 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n433), .ZN(
        u5_mult_82_ab_9__7_) );
  NOR2_X1 u5_mult_82_U482 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n431), .ZN(
        u5_mult_82_ab_9__8_) );
  NOR2_X1 u5_mult_82_U481 ( .A1(u5_mult_82_n310), .A2(u5_mult_82_n429), .ZN(
        u5_mult_82_ab_9__9_) );
  INV_X4 u5_mult_82_U479 ( .A(u6_N0), .ZN(u5_mult_82_n480) );
  INV_X4 u5_mult_82_U478 ( .A(u6_N2), .ZN(u5_mult_82_n479) );
  INV_X4 u5_mult_82_U477 ( .A(u6_N3), .ZN(u5_mult_82_n478) );
  INV_X4 u5_mult_82_U476 ( .A(u6_N10), .ZN(u5_mult_82_n477) );
  INV_X4 u5_mult_82_U475 ( .A(u6_N18), .ZN(u5_mult_82_n476) );
  INV_X4 u5_mult_82_U474 ( .A(u6_N20), .ZN(u5_mult_82_n475) );
  INV_X4 u5_mult_82_U473 ( .A(u6_N36), .ZN(u5_mult_82_n474) );
  INV_X4 u5_mult_82_U472 ( .A(fracta_mul[7]), .ZN(u5_mult_82_n473) );
  INV_X4 u5_mult_82_U471 ( .A(fracta_mul[8]), .ZN(u5_mult_82_n472) );
  INV_X4 u5_mult_82_U470 ( .A(fracta_mul[10]), .ZN(u5_mult_82_n471) );
  INV_X4 u5_mult_82_U469 ( .A(fracta_mul[11]), .ZN(u5_mult_82_n470) );
  INV_X4 u5_mult_82_U468 ( .A(fracta_mul[14]), .ZN(u5_mult_82_n469) );
  INV_X4 u5_mult_82_U467 ( .A(fracta_mul[15]), .ZN(u5_mult_82_n468) );
  INV_X4 u5_mult_82_U466 ( .A(fracta_mul[16]), .ZN(u5_mult_82_n467) );
  INV_X4 u5_mult_82_U465 ( .A(fracta_mul[17]), .ZN(u5_mult_82_n466) );
  INV_X4 u5_mult_82_U464 ( .A(fracta_mul[18]), .ZN(u5_mult_82_n465) );
  INV_X4 u5_mult_82_U463 ( .A(fracta_mul[20]), .ZN(u5_mult_82_n464) );
  INV_X4 u5_mult_82_U462 ( .A(fracta_mul[21]), .ZN(u5_mult_82_n463) );
  INV_X4 u5_mult_82_U461 ( .A(fracta_mul[25]), .ZN(u5_mult_82_n462) );
  INV_X4 u5_mult_82_U460 ( .A(fracta_mul[27]), .ZN(u5_mult_82_n461) );
  INV_X4 u5_mult_82_U459 ( .A(fracta_mul[30]), .ZN(u5_mult_82_n460) );
  INV_X4 u5_mult_82_U458 ( .A(fracta_mul[31]), .ZN(u5_mult_82_n459) );
  INV_X4 u5_mult_82_U457 ( .A(fracta_mul[32]), .ZN(u5_mult_82_n458) );
  INV_X4 u5_mult_82_U456 ( .A(fracta_mul[33]), .ZN(u5_mult_82_n457) );
  INV_X4 u5_mult_82_U455 ( .A(fracta_mul[34]), .ZN(u5_mult_82_n456) );
  INV_X4 u5_mult_82_U454 ( .A(fracta_mul[39]), .ZN(u5_mult_82_n455) );
  INV_X4 u5_mult_82_U453 ( .A(fracta_mul[43]), .ZN(u5_mult_82_n454) );
  INV_X4 u5_mult_82_U452 ( .A(fracta_mul[44]), .ZN(u5_mult_82_n453) );
  INV_X4 u5_mult_82_U451 ( .A(fracta_mul[45]), .ZN(u5_mult_82_n452) );
  INV_X4 u5_mult_82_U450 ( .A(fracta_mul[46]), .ZN(u5_mult_82_n451) );
  INV_X4 u5_mult_82_U449 ( .A(fracta_mul[50]), .ZN(u5_mult_82_n450) );
  XOR2_X2 u5_mult_82_U448 ( .A(u5_mult_82_ab_1__0_), .B(u5_mult_82_ab_0__1_), 
        .Z(u5_N1) );
  INV_X4 u5_mult_82_U447 ( .A(fracta_mul[49]), .ZN(u5_mult_82_n216) );
  INV_X4 u5_mult_82_U446 ( .A(fracta_mul[49]), .ZN(u5_mult_82_n217) );
  INV_X4 u5_mult_82_U445 ( .A(fracta_mul[48]), .ZN(u5_mult_82_n219) );
  INV_X4 u5_mult_82_U444 ( .A(fracta_mul[48]), .ZN(u5_mult_82_n220) );
  INV_X4 u5_mult_82_U443 ( .A(fracta_mul[47]), .ZN(u5_mult_82_n222) );
  INV_X4 u5_mult_82_U442 ( .A(fracta_mul[47]), .ZN(u5_mult_82_n223) );
  INV_X4 u5_mult_82_U441 ( .A(fracta_mul[51]), .ZN(u5_mult_82_n211) );
  INV_X4 u5_mult_82_U440 ( .A(n4602), .ZN(u5_mult_82_n447) );
  INV_X4 u5_mult_82_U439 ( .A(fracta_mul[44]), .ZN(u5_mult_82_n229) );
  INV_X4 u5_mult_82_U438 ( .A(fracta_mul[44]), .ZN(u5_mult_82_n230) );
  INV_X4 u5_mult_82_U437 ( .A(fracta_mul[42]), .ZN(u5_mult_82_n236) );
  INV_X4 u5_mult_82_U436 ( .A(fracta_mul[42]), .ZN(u5_mult_82_n237) );
  INV_X4 u5_mult_82_U435 ( .A(fracta_mul[42]), .ZN(u5_mult_82_n238) );
  INV_X4 u5_mult_82_U434 ( .A(u5_mult_82_n235), .ZN(u5_mult_82_n232) );
  INV_X4 u5_mult_82_U433 ( .A(u5_mult_82_n235), .ZN(u5_mult_82_n233) );
  INV_X4 u5_mult_82_U432 ( .A(fracta_mul[40]), .ZN(u5_mult_82_n244) );
  INV_X4 u5_mult_82_U431 ( .A(fracta_mul[40]), .ZN(u5_mult_82_n245) );
  INV_X4 u5_mult_82_U430 ( .A(fracta_mul[40]), .ZN(u5_mult_82_n246) );
  INV_X4 u5_mult_82_U429 ( .A(fracta_mul[45]), .ZN(u5_mult_82_n226) );
  INV_X4 u5_mult_82_U428 ( .A(fracta_mul[45]), .ZN(u5_mult_82_n227) );
  INV_X4 u5_mult_82_U427 ( .A(fracta_mul[45]), .ZN(u5_mult_82_n228) );
  INV_X4 u5_mult_82_U426 ( .A(fracta_mul[38]), .ZN(u5_mult_82_n250) );
  INV_X4 u5_mult_82_U425 ( .A(fracta_mul[38]), .ZN(u5_mult_82_n249) );
  INV_X4 u5_mult_82_U424 ( .A(fracta_mul[38]), .ZN(u5_mult_82_n251) );
  INV_X4 u5_mult_82_U423 ( .A(fracta_mul[36]), .ZN(u5_mult_82_n256) );
  INV_X4 u5_mult_82_U422 ( .A(fracta_mul[36]), .ZN(u5_mult_82_n257) );
  INV_X4 u5_mult_82_U421 ( .A(fracta_mul[37]), .ZN(u5_mult_82_n254) );
  INV_X4 u5_mult_82_U420 ( .A(fracta_mul[37]), .ZN(u5_mult_82_n255) );
  INV_X4 u5_mult_82_U419 ( .A(fracta_mul[37]), .ZN(u5_mult_82_n253) );
  INV_X4 u5_mult_82_U418 ( .A(fracta_mul[33]), .ZN(u5_mult_82_n264) );
  INV_X4 u5_mult_82_U417 ( .A(fracta_mul[33]), .ZN(u5_mult_82_n265) );
  INV_X4 u5_mult_82_U416 ( .A(fracta_mul[34]), .ZN(u5_mult_82_n262) );
  INV_X4 u5_mult_82_U415 ( .A(fracta_mul[34]), .ZN(u5_mult_82_n263) );
  INV_X4 u5_mult_82_U414 ( .A(fracta_mul[31]), .ZN(u5_mult_82_n268) );
  INV_X4 u5_mult_82_U413 ( .A(fracta_mul[32]), .ZN(u5_mult_82_n266) );
  INV_X4 u5_mult_82_U412 ( .A(fracta_mul[27]), .ZN(u5_mult_82_n279) );
  INV_X4 u5_mult_82_U411 ( .A(fracta_mul[28]), .ZN(u5_mult_82_n276) );
  INV_X4 u5_mult_82_U410 ( .A(fracta_mul[21]), .ZN(u5_mult_82_n291) );
  INV_X4 u5_mult_82_U409 ( .A(fracta_mul[22]), .ZN(u5_mult_82_n289) );
  INV_X4 u5_mult_82_U408 ( .A(fracta_mul[18]), .ZN(u5_mult_82_n295) );
  INV_X4 u5_mult_82_U407 ( .A(fracta_mul[24]), .ZN(u5_mult_82_n285) );
  INV_X4 u5_mult_82_U406 ( .A(fracta_mul[19]), .ZN(u5_mult_82_n294) );
  INV_X4 u5_mult_82_U405 ( .A(fracta_mul[23]), .ZN(u5_mult_82_n287) );
  AND2_X4 u5_mult_82_U404 ( .A1(u5_mult_82_SUMB_52__51_), .A2(
        u5_mult_82_CARRYB_52__50_), .ZN(u5_mult_82_n209) );
  AND2_X4 u5_mult_82_U403 ( .A1(u5_mult_82_ab_52__52_), .A2(
        u5_mult_82_CARRYB_52__51_), .ZN(u5_mult_82_n208) );
  INV_X4 u5_mult_82_U402 ( .A(fracta_mul[15]), .ZN(u5_mult_82_n301) );
  INV_X4 u5_mult_82_U401 ( .A(fracta_mul[16]), .ZN(u5_mult_82_n299) );
  INV_X4 u5_mult_82_U400 ( .A(fracta_mul[12]), .ZN(u5_mult_82_n306) );
  INV_X4 u5_mult_82_U399 ( .A(fracta_mul[17]), .ZN(u5_mult_82_n297) );
  XOR2_X2 u5_mult_82_U398 ( .A(u5_mult_82_CARRYB_52__0_), .B(
        u5_mult_82_SUMB_52__1_), .Z(u5_N53) );
  AND2_X4 u5_mult_82_U397 ( .A1(u5_mult_82_SUMB_52__49_), .A2(
        u5_mult_82_CARRYB_52__48_), .ZN(u5_mult_82_n206) );
  AND2_X4 u5_mult_82_U396 ( .A1(u5_mult_82_SUMB_52__47_), .A2(
        u5_mult_82_CARRYB_52__46_), .ZN(u5_mult_82_n205) );
  AND2_X4 u5_mult_82_U395 ( .A1(u5_mult_82_SUMB_52__44_), .A2(
        u5_mult_82_CARRYB_52__43_), .ZN(u5_mult_82_n204) );
  AND2_X4 u5_mult_82_U394 ( .A1(u5_mult_82_SUMB_52__42_), .A2(
        u5_mult_82_CARRYB_52__41_), .ZN(u5_mult_82_n203) );
  AND2_X4 u5_mult_82_U393 ( .A1(u5_mult_82_SUMB_52__40_), .A2(
        u5_mult_82_CARRYB_52__39_), .ZN(u5_mult_82_n202) );
  AND2_X4 u5_mult_82_U392 ( .A1(u5_mult_82_SUMB_52__45_), .A2(
        u5_mult_82_CARRYB_52__44_), .ZN(u5_mult_82_n201) );
  AND2_X4 u5_mult_82_U391 ( .A1(u5_mult_82_SUMB_52__46_), .A2(
        u5_mult_82_CARRYB_52__45_), .ZN(u5_mult_82_n200) );
  AND2_X4 u5_mult_82_U390 ( .A1(u5_mult_82_SUMB_52__41_), .A2(
        u5_mult_82_CARRYB_52__40_), .ZN(u5_mult_82_n199) );
  AND2_X4 u5_mult_82_U389 ( .A1(u5_mult_82_SUMB_52__43_), .A2(
        u5_mult_82_CARRYB_52__42_), .ZN(u5_mult_82_n198) );
  AND2_X4 u5_mult_82_U388 ( .A1(u5_mult_82_SUMB_52__48_), .A2(
        u5_mult_82_CARRYB_52__47_), .ZN(u5_mult_82_n197) );
  AND2_X4 u5_mult_82_U387 ( .A1(u5_mult_82_SUMB_52__50_), .A2(
        u5_mult_82_CARRYB_52__49_), .ZN(u5_mult_82_n196) );
  INV_X4 u5_mult_82_U386 ( .A(fracta_mul[8]), .ZN(u5_mult_82_n312) );
  INV_X4 u5_mult_82_U385 ( .A(fracta_mul[8]), .ZN(u5_mult_82_n313) );
  INV_X4 u5_mult_82_U384 ( .A(fracta_mul[7]), .ZN(u5_mult_82_n314) );
  INV_X4 u5_mult_82_U383 ( .A(fracta_mul[10]), .ZN(u5_mult_82_n309) );
  INV_X4 u5_mult_82_U382 ( .A(fracta_mul[11]), .ZN(u5_mult_82_n308) );
  INV_X4 u5_mult_82_U381 ( .A(u6_N18), .ZN(u5_mult_82_n407) );
  INV_X4 u5_mult_82_U380 ( .A(u6_N1), .ZN(u5_mult_82_n444) );
  INV_X4 u5_mult_82_U379 ( .A(fracta_mul[9]), .ZN(u5_mult_82_n310) );
  AND2_X4 u5_mult_82_U378 ( .A1(u5_mult_82_SUMB_52__36_), .A2(
        u5_mult_82_CARRYB_52__35_), .ZN(u5_mult_82_n195) );
  AND2_X4 u5_mult_82_U377 ( .A1(u5_mult_82_SUMB_52__34_), .A2(
        u5_mult_82_CARRYB_52__33_), .ZN(u5_mult_82_n194) );
  AND2_X4 u5_mult_82_U376 ( .A1(u5_mult_82_SUMB_52__33_), .A2(
        u5_mult_82_CARRYB_52__32_), .ZN(u5_mult_82_n193) );
  AND2_X4 u5_mult_82_U375 ( .A1(u5_mult_82_SUMB_52__32_), .A2(
        u5_mult_82_CARRYB_52__31_), .ZN(u5_mult_82_n192) );
  AND2_X4 u5_mult_82_U374 ( .A1(u5_mult_82_SUMB_52__30_), .A2(
        u5_mult_82_CARRYB_52__29_), .ZN(u5_mult_82_n191) );
  AND2_X4 u5_mult_82_U373 ( .A1(u5_mult_82_SUMB_52__29_), .A2(
        u5_mult_82_CARRYB_52__28_), .ZN(u5_mult_82_n190) );
  AND2_X4 u5_mult_82_U372 ( .A1(u5_mult_82_SUMB_52__20_), .A2(
        u5_mult_82_CARRYB_52__19_), .ZN(u5_mult_82_n189) );
  AND2_X4 u5_mult_82_U371 ( .A1(u5_mult_82_SUMB_52__18_), .A2(
        u5_mult_82_CARRYB_52__17_), .ZN(u5_mult_82_n188) );
  AND2_X4 u5_mult_82_U370 ( .A1(u5_mult_82_SUMB_52__17_), .A2(
        u5_mult_82_CARRYB_52__16_), .ZN(u5_mult_82_n187) );
  AND2_X4 u5_mult_82_U369 ( .A1(u5_mult_82_SUMB_52__16_), .A2(
        u5_mult_82_CARRYB_52__15_), .ZN(u5_mult_82_n186) );
  AND2_X4 u5_mult_82_U368 ( .A1(u5_mult_82_SUMB_52__24_), .A2(
        u5_mult_82_CARRYB_52__23_), .ZN(u5_mult_82_n185) );
  AND2_X4 u5_mult_82_U367 ( .A1(u5_mult_82_SUMB_52__22_), .A2(
        u5_mult_82_CARRYB_52__21_), .ZN(u5_mult_82_n184) );
  AND2_X4 u5_mult_82_U366 ( .A1(u5_mult_82_SUMB_52__21_), .A2(
        u5_mult_82_CARRYB_52__20_), .ZN(u5_mult_82_n183) );
  AND2_X4 u5_mult_82_U365 ( .A1(u5_mult_82_SUMB_52__25_), .A2(
        u5_mult_82_CARRYB_52__24_), .ZN(u5_mult_82_n182) );
  AND2_X4 u5_mult_82_U364 ( .A1(u5_mult_82_SUMB_52__27_), .A2(
        u5_mult_82_CARRYB_52__26_), .ZN(u5_mult_82_n181) );
  AND2_X4 u5_mult_82_U363 ( .A1(u5_mult_82_SUMB_52__39_), .A2(
        u5_mult_82_CARRYB_52__38_), .ZN(u5_mult_82_n180) );
  AND2_X4 u5_mult_82_U362 ( .A1(u5_mult_82_SUMB_52__38_), .A2(
        u5_mult_82_CARRYB_52__37_), .ZN(u5_mult_82_n179) );
  AND2_X4 u5_mult_82_U361 ( .A1(u5_mult_82_SUMB_52__37_), .A2(
        u5_mult_82_CARRYB_52__36_), .ZN(u5_mult_82_n178) );
  AND2_X4 u5_mult_82_U360 ( .A1(u5_mult_82_SUMB_52__35_), .A2(
        u5_mult_82_CARRYB_52__34_), .ZN(u5_mult_82_n177) );
  AND2_X4 u5_mult_82_U359 ( .A1(u5_mult_82_SUMB_52__28_), .A2(
        u5_mult_82_CARRYB_52__27_), .ZN(u5_mult_82_n176) );
  AND2_X4 u5_mult_82_U358 ( .A1(u5_mult_82_SUMB_52__26_), .A2(
        u5_mult_82_CARRYB_52__25_), .ZN(u5_mult_82_n175) );
  AND2_X4 u5_mult_82_U357 ( .A1(u5_mult_82_SUMB_52__23_), .A2(
        u5_mult_82_CARRYB_52__22_), .ZN(u5_mult_82_n174) );
  AND2_X4 u5_mult_82_U356 ( .A1(u5_mult_82_SUMB_52__31_), .A2(
        u5_mult_82_CARRYB_52__30_), .ZN(u5_mult_82_n173) );
  AND2_X4 u5_mult_82_U355 ( .A1(u5_mult_82_SUMB_52__19_), .A2(
        u5_mult_82_CARRYB_52__18_), .ZN(u5_mult_82_n172) );
  INV_X4 u5_mult_82_U354 ( .A(fracta_mul[6]), .ZN(u5_mult_82_n318) );
  XOR2_X2 u5_mult_82_U353 ( .A(u5_mult_82_ab_1__1_), .B(u5_mult_82_ab_0__2_), 
        .Z(u5_mult_82_n171) );
  INV_X4 u5_mult_82_U352 ( .A(fracta_mul[0]), .ZN(u5_mult_82_n333) );
  INV_X4 u5_mult_82_U351 ( .A(fracta_mul[0]), .ZN(u5_mult_82_n334) );
  INV_X4 u5_mult_82_U350 ( .A(fracta_mul[0]), .ZN(u5_mult_82_n335) );
  INV_X4 u5_mult_82_U349 ( .A(fracta_mul[3]), .ZN(u5_mult_82_n325) );
  INV_X4 u5_mult_82_U348 ( .A(fracta_mul[3]), .ZN(u5_mult_82_n326) );
  INV_X4 u5_mult_82_U347 ( .A(fracta_mul[4]), .ZN(u5_mult_82_n323) );
  INV_X4 u5_mult_82_U346 ( .A(fracta_mul[4]), .ZN(u5_mult_82_n324) );
  INV_X4 u5_mult_82_U345 ( .A(fracta_mul[1]), .ZN(u5_mult_82_n331) );
  INV_X4 u5_mult_82_U344 ( .A(fracta_mul[1]), .ZN(u5_mult_82_n332) );
  INV_X4 u5_mult_82_U343 ( .A(fracta_mul[5]), .ZN(u5_mult_82_n320) );
  INV_X4 u5_mult_82_U342 ( .A(fracta_mul[5]), .ZN(u5_mult_82_n321) );
  INV_X4 u5_mult_82_U341 ( .A(fracta_mul[5]), .ZN(u5_mult_82_n322) );
  INV_X4 u5_mult_82_U340 ( .A(fracta_mul[2]), .ZN(u5_mult_82_n328) );
  INV_X4 u5_mult_82_U339 ( .A(fracta_mul[2]), .ZN(u5_mult_82_n329) );
  INV_X4 u5_mult_82_U338 ( .A(u6_N43), .ZN(u5_mult_82_n357) );
  INV_X4 u5_mult_82_U337 ( .A(u6_N49), .ZN(u5_mult_82_n344) );
  INV_X4 u5_mult_82_U336 ( .A(u6_N19), .ZN(u5_mult_82_n405) );
  INV_X4 u5_mult_82_U335 ( .A(u6_N15), .ZN(u5_mult_82_n414) );
  INV_X4 u5_mult_82_U334 ( .A(u6_N15), .ZN(u5_mult_82_n415) );
  INV_X4 u5_mult_82_U333 ( .A(u6_N16), .ZN(u5_mult_82_n411) );
  INV_X4 u5_mult_82_U332 ( .A(u6_N16), .ZN(u5_mult_82_n412) );
  INV_X4 u5_mult_82_U331 ( .A(u6_N12), .ZN(u5_mult_82_n423) );
  INV_X4 u5_mult_82_U330 ( .A(u6_N12), .ZN(u5_mult_82_n424) );
  INV_X4 u5_mult_82_U329 ( .A(u6_N13), .ZN(u5_mult_82_n420) );
  INV_X4 u5_mult_82_U328 ( .A(u6_N13), .ZN(u5_mult_82_n421) );
  INV_X4 u5_mult_82_U327 ( .A(u6_N14), .ZN(u5_mult_82_n417) );
  INV_X4 u5_mult_82_U326 ( .A(u6_N14), .ZN(u5_mult_82_n418) );
  AND2_X4 u5_mult_82_U325 ( .A1(u5_mult_82_SUMB_52__14_), .A2(
        u5_mult_82_CARRYB_52__13_), .ZN(u5_mult_82_n170) );
  AND2_X4 u5_mult_82_U324 ( .A1(u5_mult_82_SUMB_52__13_), .A2(
        u5_mult_82_CARRYB_52__12_), .ZN(u5_mult_82_n169) );
  AND2_X4 u5_mult_82_U323 ( .A1(u5_mult_82_SUMB_52__15_), .A2(
        u5_mult_82_CARRYB_52__14_), .ZN(u5_mult_82_n168) );
  AND2_X4 u5_mult_82_U322 ( .A1(u5_mult_82_SUMB_52__11_), .A2(
        u5_mult_82_CARRYB_52__10_), .ZN(u5_mult_82_n167) );
  AND2_X4 u5_mult_82_U321 ( .A1(u5_mult_82_SUMB_52__9_), .A2(
        u5_mult_82_CARRYB_52__8_), .ZN(u5_mult_82_n166) );
  AND2_X4 u5_mult_82_U320 ( .A1(u5_mult_82_SUMB_52__8_), .A2(
        u5_mult_82_CARRYB_52__7_), .ZN(u5_mult_82_n165) );
  AND2_X4 u5_mult_82_U319 ( .A1(u5_mult_82_SUMB_52__6_), .A2(
        u5_mult_82_CARRYB_52__5_), .ZN(u5_mult_82_n164) );
  AND2_X4 u5_mult_82_U318 ( .A1(u5_mult_82_SUMB_52__4_), .A2(
        u5_mult_82_CARRYB_52__3_), .ZN(u5_mult_82_n163) );
  AND2_X4 u5_mult_82_U317 ( .A1(u5_mult_82_SUMB_52__12_), .A2(
        u5_mult_82_CARRYB_52__11_), .ZN(u5_mult_82_n162) );
  AND2_X4 u5_mult_82_U316 ( .A1(u5_mult_82_SUMB_52__10_), .A2(
        u5_mult_82_CARRYB_52__9_), .ZN(u5_mult_82_n161) );
  AND2_X4 u5_mult_82_U315 ( .A1(u5_mult_82_SUMB_52__7_), .A2(
        u5_mult_82_CARRYB_52__6_), .ZN(u5_mult_82_n160) );
  AND2_X4 u5_mult_82_U314 ( .A1(u5_mult_82_SUMB_52__5_), .A2(
        u5_mult_82_CARRYB_52__4_), .ZN(u5_mult_82_n159) );
  INV_X4 u5_mult_82_U313 ( .A(u6_N50), .ZN(u5_mult_82_n342) );
  XOR2_X2 u5_mult_82_U312 ( .A(u5_mult_82_ab_1__2_), .B(u5_mult_82_ab_0__3_), 
        .Z(u5_mult_82_n158) );
  XOR2_X2 u5_mult_82_U311 ( .A(u5_mult_82_ab_1__3_), .B(u5_mult_82_ab_0__4_), 
        .Z(u5_mult_82_n157) );
  XOR2_X2 u5_mult_82_U310 ( .A(u5_mult_82_ab_1__4_), .B(u5_mult_82_ab_0__5_), 
        .Z(u5_mult_82_n156) );
  XOR2_X2 u5_mult_82_U309 ( .A(u5_mult_82_ab_1__5_), .B(u5_mult_82_ab_0__6_), 
        .Z(u5_mult_82_n155) );
  XOR2_X2 u5_mult_82_U308 ( .A(u5_mult_82_ab_1__6_), .B(u5_mult_82_ab_0__7_), 
        .Z(u5_mult_82_n154) );
  XOR2_X2 u5_mult_82_U307 ( .A(u5_mult_82_ab_1__7_), .B(u5_mult_82_ab_0__8_), 
        .Z(u5_mult_82_n153) );
  XOR2_X2 u5_mult_82_U306 ( .A(u5_mult_82_ab_1__8_), .B(u5_mult_82_ab_0__9_), 
        .Z(u5_mult_82_n152) );
  XOR2_X2 u5_mult_82_U305 ( .A(u5_mult_82_ab_1__9_), .B(u5_mult_82_ab_0__10_), 
        .Z(u5_mult_82_n151) );
  XOR2_X2 u5_mult_82_U304 ( .A(u5_mult_82_ab_1__10_), .B(u5_mult_82_ab_0__11_), 
        .Z(u5_mult_82_n150) );
  XOR2_X2 u5_mult_82_U303 ( .A(u5_mult_82_ab_1__11_), .B(u5_mult_82_ab_0__12_), 
        .Z(u5_mult_82_n149) );
  XOR2_X2 u5_mult_82_U302 ( .A(u5_mult_82_ab_1__12_), .B(u5_mult_82_ab_0__13_), 
        .Z(u5_mult_82_n148) );
  XOR2_X2 u5_mult_82_U301 ( .A(u5_mult_82_ab_1__13_), .B(u5_mult_82_ab_0__14_), 
        .Z(u5_mult_82_n147) );
  XOR2_X2 u5_mult_82_U300 ( .A(u5_mult_82_ab_1__14_), .B(u5_mult_82_ab_0__15_), 
        .Z(u5_mult_82_n146) );
  XOR2_X2 u5_mult_82_U299 ( .A(u5_mult_82_ab_1__15_), .B(u5_mult_82_ab_0__16_), 
        .Z(u5_mult_82_n145) );
  XOR2_X2 u5_mult_82_U298 ( .A(u5_mult_82_ab_1__16_), .B(u5_mult_82_ab_0__17_), 
        .Z(u5_mult_82_n144) );
  XOR2_X2 u5_mult_82_U297 ( .A(u5_mult_82_ab_1__17_), .B(u5_mult_82_ab_0__18_), 
        .Z(u5_mult_82_n143) );
  XOR2_X2 u5_mult_82_U296 ( .A(u5_mult_82_ab_1__18_), .B(u5_mult_82_ab_0__19_), 
        .Z(u5_mult_82_n142) );
  XOR2_X2 u5_mult_82_U295 ( .A(u5_mult_82_ab_1__19_), .B(u5_mult_82_ab_0__20_), 
        .Z(u5_mult_82_n141) );
  XOR2_X2 u5_mult_82_U294 ( .A(u5_mult_82_ab_1__20_), .B(u5_mult_82_ab_0__21_), 
        .Z(u5_mult_82_n140) );
  XOR2_X2 u5_mult_82_U293 ( .A(u5_mult_82_ab_1__21_), .B(u5_mult_82_ab_0__22_), 
        .Z(u5_mult_82_n139) );
  XOR2_X2 u5_mult_82_U292 ( .A(u5_mult_82_ab_1__22_), .B(u5_mult_82_ab_0__23_), 
        .Z(u5_mult_82_n138) );
  XOR2_X2 u5_mult_82_U291 ( .A(u5_mult_82_ab_1__23_), .B(u5_mult_82_ab_0__24_), 
        .Z(u5_mult_82_n137) );
  XOR2_X2 u5_mult_82_U290 ( .A(u5_mult_82_ab_1__24_), .B(u5_mult_82_ab_0__25_), 
        .Z(u5_mult_82_n136) );
  XOR2_X2 u5_mult_82_U289 ( .A(u5_mult_82_ab_1__25_), .B(u5_mult_82_ab_0__26_), 
        .Z(u5_mult_82_n135) );
  XOR2_X2 u5_mult_82_U288 ( .A(u5_mult_82_ab_1__26_), .B(u5_mult_82_ab_0__27_), 
        .Z(u5_mult_82_n134) );
  XOR2_X2 u5_mult_82_U287 ( .A(u5_mult_82_ab_1__27_), .B(u5_mult_82_ab_0__28_), 
        .Z(u5_mult_82_n133) );
  XOR2_X2 u5_mult_82_U286 ( .A(u5_mult_82_ab_1__28_), .B(u5_mult_82_ab_0__29_), 
        .Z(u5_mult_82_n132) );
  XOR2_X2 u5_mult_82_U285 ( .A(u5_mult_82_ab_1__29_), .B(u5_mult_82_ab_0__30_), 
        .Z(u5_mult_82_n131) );
  XOR2_X2 u5_mult_82_U284 ( .A(u5_mult_82_ab_1__30_), .B(u5_mult_82_ab_0__31_), 
        .Z(u5_mult_82_n130) );
  XOR2_X2 u5_mult_82_U283 ( .A(u5_mult_82_ab_1__31_), .B(u5_mult_82_ab_0__32_), 
        .Z(u5_mult_82_n129) );
  XOR2_X2 u5_mult_82_U282 ( .A(u5_mult_82_ab_1__32_), .B(u5_mult_82_ab_0__33_), 
        .Z(u5_mult_82_n128) );
  XOR2_X2 u5_mult_82_U281 ( .A(u5_mult_82_ab_1__33_), .B(u5_mult_82_ab_0__34_), 
        .Z(u5_mult_82_n127) );
  XOR2_X2 u5_mult_82_U280 ( .A(u5_mult_82_ab_1__34_), .B(u5_mult_82_ab_0__35_), 
        .Z(u5_mult_82_n126) );
  XOR2_X2 u5_mult_82_U279 ( .A(u5_mult_82_ab_1__35_), .B(u5_mult_82_ab_0__36_), 
        .Z(u5_mult_82_n125) );
  XOR2_X2 u5_mult_82_U278 ( .A(u5_mult_82_ab_1__36_), .B(u5_mult_82_ab_0__37_), 
        .Z(u5_mult_82_n124) );
  XOR2_X2 u5_mult_82_U277 ( .A(u5_mult_82_ab_1__37_), .B(u5_mult_82_ab_0__38_), 
        .Z(u5_mult_82_n123) );
  XOR2_X2 u5_mult_82_U276 ( .A(u5_mult_82_ab_1__38_), .B(u5_mult_82_ab_0__39_), 
        .Z(u5_mult_82_n122) );
  XOR2_X2 u5_mult_82_U275 ( .A(u5_mult_82_ab_1__39_), .B(u5_mult_82_ab_0__40_), 
        .Z(u5_mult_82_n121) );
  XOR2_X2 u5_mult_82_U274 ( .A(u5_mult_82_ab_1__40_), .B(u5_mult_82_ab_0__41_), 
        .Z(u5_mult_82_n120) );
  XOR2_X2 u5_mult_82_U273 ( .A(u5_mult_82_ab_1__41_), .B(u5_mult_82_ab_0__42_), 
        .Z(u5_mult_82_n119) );
  XOR2_X2 u5_mult_82_U272 ( .A(u5_mult_82_ab_1__42_), .B(u5_mult_82_ab_0__43_), 
        .Z(u5_mult_82_n118) );
  XOR2_X2 u5_mult_82_U271 ( .A(u5_mult_82_ab_1__43_), .B(u5_mult_82_ab_0__44_), 
        .Z(u5_mult_82_n117) );
  XOR2_X2 u5_mult_82_U270 ( .A(u5_mult_82_ab_1__44_), .B(u5_mult_82_ab_0__45_), 
        .Z(u5_mult_82_n116) );
  XOR2_X2 u5_mult_82_U269 ( .A(u5_mult_82_ab_1__45_), .B(u5_mult_82_ab_0__46_), 
        .Z(u5_mult_82_n115) );
  XOR2_X2 u5_mult_82_U268 ( .A(u5_mult_82_ab_1__46_), .B(u5_mult_82_ab_0__47_), 
        .Z(u5_mult_82_n114) );
  XOR2_X2 u5_mult_82_U267 ( .A(u5_mult_82_ab_1__47_), .B(u5_mult_82_ab_0__48_), 
        .Z(u5_mult_82_n113) );
  XOR2_X2 u5_mult_82_U266 ( .A(u5_mult_82_ab_1__48_), .B(u5_mult_82_ab_0__49_), 
        .Z(u5_mult_82_n112) );
  XOR2_X2 u5_mult_82_U265 ( .A(u5_mult_82_ab_1__49_), .B(u5_mult_82_ab_0__50_), 
        .Z(u5_mult_82_n111) );
  XOR2_X2 u5_mult_82_U264 ( .A(u5_mult_82_ab_1__50_), .B(u5_mult_82_ab_0__51_), 
        .Z(u5_mult_82_n110) );
  AND2_X4 u5_mult_82_U263 ( .A1(u5_mult_82_ab_0__51_), .A2(
        u5_mult_82_ab_1__50_), .ZN(u5_mult_82_n109) );
  AND2_X4 u5_mult_82_U262 ( .A1(u5_mult_82_SUMB_52__3_), .A2(
        u5_mult_82_CARRYB_52__2_), .ZN(u5_mult_82_n108) );
  AND2_X4 u5_mult_82_U261 ( .A1(u5_mult_82_SUMB_52__1_), .A2(
        u5_mult_82_CARRYB_52__0_), .ZN(u5_mult_82_n107) );
  AND2_X4 u5_mult_82_U260 ( .A1(u5_mult_82_SUMB_52__2_), .A2(
        u5_mult_82_CARRYB_52__1_), .ZN(u5_mult_82_n106) );
  AND2_X4 u5_mult_82_U259 ( .A1(u5_mult_82_ab_0__52_), .A2(
        u5_mult_82_ab_1__51_), .ZN(u5_mult_82_n105) );
  INV_X4 u5_mult_82_U258 ( .A(n4602), .ZN(u5_mult_82_n448) );
  INV_X4 u5_mult_82_U257 ( .A(fracta_mul[50]), .ZN(u5_mult_82_n213) );
  INV_X4 u5_mult_82_U256 ( .A(fracta_mul[46]), .ZN(u5_mult_82_n225) );
  INV_X4 u5_mult_82_U255 ( .A(fracta_mul[51]), .ZN(u5_mult_82_n212) );
  INV_X4 u5_mult_82_U254 ( .A(fracta_mul[49]), .ZN(u5_mult_82_n215) );
  INV_X4 u5_mult_82_U253 ( .A(fracta_mul[48]), .ZN(u5_mult_82_n218) );
  INV_X4 u5_mult_82_U252 ( .A(fracta_mul[47]), .ZN(u5_mult_82_n221) );
  INV_X4 u5_mult_82_U251 ( .A(fracta_mul[44]), .ZN(u5_mult_82_n231) );
  INV_X4 u5_mult_82_U250 ( .A(fracta_mul[42]), .ZN(u5_mult_82_n239) );
  INV_X4 u5_mult_82_U249 ( .A(u5_mult_82_n235), .ZN(u5_mult_82_n234) );
  INV_X4 u5_mult_82_U248 ( .A(fracta_mul[41]), .ZN(u5_mult_82_n240) );
  INV_X4 u5_mult_82_U247 ( .A(fracta_mul[41]), .ZN(u5_mult_82_n241) );
  INV_X4 u5_mult_82_U246 ( .A(fracta_mul[41]), .ZN(u5_mult_82_n242) );
  INV_X4 u5_mult_82_U245 ( .A(fracta_mul[39]), .ZN(u5_mult_82_n247) );
  INV_X4 u5_mult_82_U244 ( .A(fracta_mul[38]), .ZN(u5_mult_82_n252) );
  INV_X4 u5_mult_82_U243 ( .A(fracta_mul[35]), .ZN(u5_mult_82_n259) );
  INV_X4 u5_mult_82_U242 ( .A(fracta_mul[35]), .ZN(u5_mult_82_n260) );
  INV_X4 u5_mult_82_U241 ( .A(fracta_mul[36]), .ZN(u5_mult_82_n258) );
  INV_X4 u5_mult_82_U240 ( .A(fracta_mul[25]), .ZN(u5_mult_82_n283) );
  INV_X4 u5_mult_82_U239 ( .A(fracta_mul[30]), .ZN(u5_mult_82_n270) );
  INV_X4 u5_mult_82_U238 ( .A(fracta_mul[30]), .ZN(u5_mult_82_n271) );
  INV_X4 u5_mult_82_U237 ( .A(fracta_mul[29]), .ZN(u5_mult_82_n273) );
  INV_X4 u5_mult_82_U236 ( .A(fracta_mul[29]), .ZN(u5_mult_82_n272) );
  INV_X4 u5_mult_82_U235 ( .A(fracta_mul[27]), .ZN(u5_mult_82_n278) );
  INV_X4 u5_mult_82_U234 ( .A(fracta_mul[32]), .ZN(u5_mult_82_n267) );
  INV_X4 u5_mult_82_U233 ( .A(fracta_mul[28]), .ZN(u5_mult_82_n275) );
  INV_X4 u5_mult_82_U232 ( .A(fracta_mul[26]), .ZN(u5_mult_82_n280) );
  INV_X4 u5_mult_82_U231 ( .A(fracta_mul[17]), .ZN(u5_mult_82_n298) );
  INV_X4 u5_mult_82_U230 ( .A(fracta_mul[13]), .ZN(u5_mult_82_n304) );
  XOR2_X2 u5_mult_82_U229 ( .A(u5_mult_82_CARRYB_52__49_), .B(
        u5_mult_82_SUMB_52__50_), .Z(u5_mult_82_n104) );
  XOR2_X2 u5_mult_82_U228 ( .A(u5_mult_82_CARRYB_52__47_), .B(
        u5_mult_82_SUMB_52__48_), .Z(u5_mult_82_n103) );
  XOR2_X2 u5_mult_82_U227 ( .A(u5_mult_82_CARRYB_52__44_), .B(
        u5_mult_82_SUMB_52__45_), .Z(u5_mult_82_n102) );
  XOR2_X2 u5_mult_82_U226 ( .A(u5_mult_82_CARRYB_52__42_), .B(
        u5_mult_82_SUMB_52__43_), .Z(u5_mult_82_n101) );
  XOR2_X2 u5_mult_82_U225 ( .A(u5_mult_82_CARRYB_52__45_), .B(
        u5_mult_82_SUMB_52__46_), .Z(u5_mult_82_n100) );
  XOR2_X2 u5_mult_82_U224 ( .A(u5_mult_82_CARRYB_52__46_), .B(
        u5_mult_82_SUMB_52__47_), .Z(u5_mult_82_n99) );
  XOR2_X2 u5_mult_82_U223 ( .A(u5_mult_82_CARRYB_52__41_), .B(
        u5_mult_82_SUMB_52__42_), .Z(u5_mult_82_n98) );
  XOR2_X2 u5_mult_82_U222 ( .A(u5_mult_82_CARRYB_52__43_), .B(
        u5_mult_82_SUMB_52__44_), .Z(u5_mult_82_n97) );
  XOR2_X2 u5_mult_82_U221 ( .A(u5_mult_82_CARRYB_52__48_), .B(
        u5_mult_82_SUMB_52__49_), .Z(u5_mult_82_n96) );
  XOR2_X2 u5_mult_82_U220 ( .A(u5_mult_82_CARRYB_52__50_), .B(
        u5_mult_82_SUMB_52__51_), .Z(u5_mult_82_n95) );
  XOR2_X2 u5_mult_82_U219 ( .A(u5_mult_82_CARRYB_52__51_), .B(
        u5_mult_82_ab_52__52_), .Z(u5_mult_82_n94) );
  INV_X4 u5_mult_82_U218 ( .A(u6_N1), .ZN(u5_mult_82_n443) );
  INV_X4 u5_mult_82_U217 ( .A(u6_N1), .ZN(u5_mult_82_n445) );
  INV_X4 u5_mult_82_U216 ( .A(u6_N3), .ZN(u5_mult_82_n441) );
  XOR2_X2 u5_mult_82_U215 ( .A(u5_mult_82_CARRYB_52__36_), .B(
        u5_mult_82_SUMB_52__37_), .Z(u5_mult_82_n93) );
  XOR2_X2 u5_mult_82_U214 ( .A(u5_mult_82_CARRYB_52__34_), .B(
        u5_mult_82_SUMB_52__35_), .Z(u5_mult_82_n92) );
  XOR2_X2 u5_mult_82_U213 ( .A(u5_mult_82_CARRYB_52__33_), .B(
        u5_mult_82_SUMB_52__34_), .Z(u5_mult_82_n91) );
  XOR2_X2 u5_mult_82_U212 ( .A(u5_mult_82_CARRYB_52__32_), .B(
        u5_mult_82_SUMB_52__33_), .Z(u5_mult_82_n90) );
  XOR2_X2 u5_mult_82_U211 ( .A(u5_mult_82_CARRYB_52__30_), .B(
        u5_mult_82_SUMB_52__31_), .Z(u5_mult_82_n89) );
  XOR2_X2 u5_mult_82_U210 ( .A(u5_mult_82_CARRYB_52__29_), .B(
        u5_mult_82_SUMB_52__30_), .Z(u5_mult_82_n88) );
  XOR2_X2 u5_mult_82_U209 ( .A(u5_mult_82_CARRYB_52__20_), .B(
        u5_mult_82_SUMB_52__21_), .Z(u5_mult_82_n87) );
  XOR2_X2 u5_mult_82_U208 ( .A(u5_mult_82_CARRYB_52__24_), .B(
        u5_mult_82_SUMB_52__25_), .Z(u5_mult_82_n86) );
  XOR2_X2 u5_mult_82_U207 ( .A(u5_mult_82_CARRYB_52__22_), .B(
        u5_mult_82_SUMB_52__23_), .Z(u5_mult_82_n85) );
  XOR2_X2 u5_mult_82_U206 ( .A(u5_mult_82_CARRYB_52__21_), .B(
        u5_mult_82_SUMB_52__22_), .Z(u5_mult_82_n84) );
  XOR2_X2 u5_mult_82_U205 ( .A(u5_mult_82_CARRYB_52__25_), .B(
        u5_mult_82_SUMB_52__26_), .Z(u5_mult_82_n83) );
  XOR2_X2 u5_mult_82_U204 ( .A(u5_mult_82_CARRYB_52__27_), .B(
        u5_mult_82_SUMB_52__28_), .Z(u5_mult_82_n82) );
  XOR2_X2 u5_mult_82_U203 ( .A(u5_mult_82_CARRYB_52__40_), .B(
        u5_mult_82_SUMB_52__41_), .Z(u5_mult_82_n81) );
  XOR2_X2 u5_mult_82_U202 ( .A(u5_mult_82_CARRYB_52__39_), .B(
        u5_mult_82_SUMB_52__40_), .Z(u5_mult_82_n80) );
  XOR2_X2 u5_mult_82_U201 ( .A(u5_mult_82_CARRYB_52__38_), .B(
        u5_mult_82_SUMB_52__39_), .Z(u5_mult_82_n79) );
  XOR2_X2 u5_mult_82_U200 ( .A(u5_mult_82_CARRYB_52__37_), .B(
        u5_mult_82_SUMB_52__38_), .Z(u5_mult_82_n78) );
  XOR2_X2 u5_mult_82_U199 ( .A(u5_mult_82_CARRYB_52__31_), .B(
        u5_mult_82_SUMB_52__32_), .Z(u5_mult_82_n77) );
  XOR2_X2 u5_mult_82_U198 ( .A(u5_mult_82_CARRYB_52__35_), .B(
        u5_mult_82_SUMB_52__36_), .Z(u5_mult_82_n76) );
  XOR2_X2 u5_mult_82_U197 ( .A(u5_mult_82_CARRYB_52__28_), .B(
        u5_mult_82_SUMB_52__29_), .Z(u5_mult_82_n75) );
  XOR2_X2 u5_mult_82_U196 ( .A(u5_mult_82_CARRYB_52__26_), .B(
        u5_mult_82_SUMB_52__27_), .Z(u5_mult_82_n74) );
  XOR2_X2 u5_mult_82_U195 ( .A(u5_mult_82_CARRYB_52__23_), .B(
        u5_mult_82_SUMB_52__24_), .Z(u5_mult_82_n73) );
  AND2_X4 u5_mult_82_U194 ( .A1(u5_mult_82_ab_0__1_), .A2(u5_mult_82_ab_1__0_), 
        .ZN(u5_mult_82_n72) );
  INV_X4 u5_mult_82_U193 ( .A(u6_N37), .ZN(u5_mult_82_n371) );
  INV_X4 u5_mult_82_U192 ( .A(u6_N30), .ZN(u5_mult_82_n384) );
  INV_X4 u5_mult_82_U191 ( .A(u6_N31), .ZN(u5_mult_82_n382) );
  INV_X4 u5_mult_82_U190 ( .A(u6_N33), .ZN(u5_mult_82_n378) );
  INV_X4 u5_mult_82_U189 ( .A(u6_N35), .ZN(u5_mult_82_n374) );
  INV_X4 u5_mult_82_U188 ( .A(u6_N39), .ZN(u5_mult_82_n366) );
  INV_X4 u5_mult_82_U187 ( .A(u6_N40), .ZN(u5_mult_82_n364) );
  INV_X4 u5_mult_82_U186 ( .A(u6_N41), .ZN(u5_mult_82_n362) );
  INV_X4 u5_mult_82_U185 ( .A(u6_N45), .ZN(u5_mult_82_n352) );
  INV_X4 u5_mult_82_U184 ( .A(u6_N46), .ZN(u5_mult_82_n350) );
  INV_X4 u5_mult_82_U183 ( .A(u6_N47), .ZN(u5_mult_82_n348) );
  INV_X4 u5_mult_82_U182 ( .A(u6_N48), .ZN(u5_mult_82_n346) );
  INV_X4 u5_mult_82_U181 ( .A(u6_N21), .ZN(u5_mult_82_n402) );
  INV_X4 u5_mult_82_U180 ( .A(u6_N34), .ZN(u5_mult_82_n376) );
  INV_X4 u5_mult_82_U179 ( .A(u6_N26), .ZN(u5_mult_82_n392) );
  INV_X4 u5_mult_82_U178 ( .A(u6_N29), .ZN(u5_mult_82_n386) );
  INV_X4 u5_mult_82_U177 ( .A(u6_N23), .ZN(u5_mult_82_n398) );
  INV_X4 u5_mult_82_U176 ( .A(u6_N24), .ZN(u5_mult_82_n396) );
  INV_X4 u5_mult_82_U175 ( .A(u6_N25), .ZN(u5_mult_82_n394) );
  INV_X4 u5_mult_82_U174 ( .A(u6_N38), .ZN(u5_mult_82_n367) );
  INV_X4 u5_mult_82_U173 ( .A(u6_N38), .ZN(u5_mult_82_n368) );
  INV_X4 u5_mult_82_U172 ( .A(u6_N42), .ZN(u5_mult_82_n359) );
  INV_X4 u5_mult_82_U171 ( .A(u6_N42), .ZN(u5_mult_82_n360) );
  INV_X4 u5_mult_82_U170 ( .A(u6_N44), .ZN(u5_mult_82_n354) );
  INV_X4 u5_mult_82_U169 ( .A(u6_N44), .ZN(u5_mult_82_n355) );
  INV_X4 u5_mult_82_U168 ( .A(u6_N22), .ZN(u5_mult_82_n400) );
  INV_X4 u5_mult_82_U167 ( .A(u6_N27), .ZN(u5_mult_82_n390) );
  INV_X4 u5_mult_82_U166 ( .A(u6_N28), .ZN(u5_mult_82_n388) );
  INV_X4 u5_mult_82_U165 ( .A(fracta_mul[2]), .ZN(u5_mult_82_n327) );
  XOR2_X2 u5_mult_82_U164 ( .A(u5_mult_82_CARRYB_52__18_), .B(
        u5_mult_82_SUMB_52__19_), .Z(u5_mult_82_n71) );
  XOR2_X2 u5_mult_82_U163 ( .A(u5_mult_82_CARRYB_52__17_), .B(
        u5_mult_82_SUMB_52__18_), .Z(u5_mult_82_n70) );
  XOR2_X2 u5_mult_82_U162 ( .A(u5_mult_82_CARRYB_52__16_), .B(
        u5_mult_82_SUMB_52__17_), .Z(u5_mult_82_n69) );
  XOR2_X2 u5_mult_82_U161 ( .A(u5_mult_82_CARRYB_52__14_), .B(
        u5_mult_82_SUMB_52__15_), .Z(u5_mult_82_n68) );
  XOR2_X2 u5_mult_82_U160 ( .A(u5_mult_82_CARRYB_52__13_), .B(
        u5_mult_82_SUMB_52__14_), .Z(u5_mult_82_n67) );
  XOR2_X2 u5_mult_82_U159 ( .A(u5_mult_82_CARRYB_52__15_), .B(
        u5_mult_82_SUMB_52__16_), .Z(u5_mult_82_n66) );
  XOR2_X2 u5_mult_82_U158 ( .A(u5_mult_82_CARRYB_52__11_), .B(
        u5_mult_82_SUMB_52__12_), .Z(u5_mult_82_n65) );
  XOR2_X2 u5_mult_82_U157 ( .A(u5_mult_82_CARRYB_52__9_), .B(
        u5_mult_82_SUMB_52__10_), .Z(u5_mult_82_n64) );
  XOR2_X2 u5_mult_82_U156 ( .A(u5_mult_82_CARRYB_52__8_), .B(
        u5_mult_82_SUMB_52__9_), .Z(u5_mult_82_n63) );
  XOR2_X2 u5_mult_82_U155 ( .A(u5_mult_82_CARRYB_52__6_), .B(
        u5_mult_82_SUMB_52__7_), .Z(u5_mult_82_n62) );
  XOR2_X2 u5_mult_82_U154 ( .A(u5_mult_82_CARRYB_52__4_), .B(
        u5_mult_82_SUMB_52__5_), .Z(u5_mult_82_n61) );
  XOR2_X2 u5_mult_82_U153 ( .A(u5_mult_82_CARRYB_52__19_), .B(
        u5_mult_82_SUMB_52__20_), .Z(u5_mult_82_n60) );
  XOR2_X2 u5_mult_82_U152 ( .A(u5_mult_82_CARRYB_52__7_), .B(
        u5_mult_82_SUMB_52__8_), .Z(u5_mult_82_n59) );
  XOR2_X2 u5_mult_82_U151 ( .A(u5_mult_82_CARRYB_52__5_), .B(
        u5_mult_82_SUMB_52__6_), .Z(u5_mult_82_n58) );
  XOR2_X2 u5_mult_82_U150 ( .A(u5_mult_82_CARRYB_52__12_), .B(
        u5_mult_82_SUMB_52__13_), .Z(u5_mult_82_n57) );
  XOR2_X2 u5_mult_82_U149 ( .A(u5_mult_82_CARRYB_52__10_), .B(
        u5_mult_82_SUMB_52__11_), .Z(u5_mult_82_n56) );
  AND2_X4 u5_mult_82_U148 ( .A1(u5_mult_82_ab_0__6_), .A2(u5_mult_82_ab_1__5_), 
        .ZN(u5_mult_82_n55) );
  AND2_X4 u5_mult_82_U147 ( .A1(u5_mult_82_ab_0__8_), .A2(u5_mult_82_ab_1__7_), 
        .ZN(u5_mult_82_n54) );
  AND2_X4 u5_mult_82_U146 ( .A1(u5_mult_82_ab_0__10_), .A2(u5_mult_82_ab_1__9_), .ZN(u5_mult_82_n53) );
  AND2_X4 u5_mult_82_U145 ( .A1(u5_mult_82_ab_0__11_), .A2(
        u5_mult_82_ab_1__10_), .ZN(u5_mult_82_n52) );
  AND2_X4 u5_mult_82_U144 ( .A1(u5_mult_82_ab_0__12_), .A2(
        u5_mult_82_ab_1__11_), .ZN(u5_mult_82_n51) );
  AND2_X4 u5_mult_82_U143 ( .A1(u5_mult_82_ab_0__13_), .A2(
        u5_mult_82_ab_1__12_), .ZN(u5_mult_82_n50) );
  AND2_X4 u5_mult_82_U142 ( .A1(u5_mult_82_ab_0__14_), .A2(
        u5_mult_82_ab_1__13_), .ZN(u5_mult_82_n49) );
  AND2_X4 u5_mult_82_U141 ( .A1(u5_mult_82_ab_0__15_), .A2(
        u5_mult_82_ab_1__14_), .ZN(u5_mult_82_n48) );
  AND2_X4 u5_mult_82_U140 ( .A1(u5_mult_82_ab_0__16_), .A2(
        u5_mult_82_ab_1__15_), .ZN(u5_mult_82_n47) );
  AND2_X4 u5_mult_82_U139 ( .A1(u5_mult_82_ab_0__17_), .A2(
        u5_mult_82_ab_1__16_), .ZN(u5_mult_82_n46) );
  AND2_X4 u5_mult_82_U138 ( .A1(u5_mult_82_ab_0__18_), .A2(
        u5_mult_82_ab_1__17_), .ZN(u5_mult_82_n45) );
  AND2_X4 u5_mult_82_U137 ( .A1(u5_mult_82_ab_0__19_), .A2(
        u5_mult_82_ab_1__18_), .ZN(u5_mult_82_n44) );
  AND2_X4 u5_mult_82_U136 ( .A1(u5_mult_82_ab_0__20_), .A2(
        u5_mult_82_ab_1__19_), .ZN(u5_mult_82_n43) );
  AND2_X4 u5_mult_82_U135 ( .A1(u5_mult_82_ab_0__21_), .A2(
        u5_mult_82_ab_1__20_), .ZN(u5_mult_82_n42) );
  AND2_X4 u5_mult_82_U134 ( .A1(u5_mult_82_ab_0__22_), .A2(
        u5_mult_82_ab_1__21_), .ZN(u5_mult_82_n41) );
  AND2_X4 u5_mult_82_U133 ( .A1(u5_mult_82_ab_0__23_), .A2(
        u5_mult_82_ab_1__22_), .ZN(u5_mult_82_n40) );
  AND2_X4 u5_mult_82_U132 ( .A1(u5_mult_82_ab_0__24_), .A2(
        u5_mult_82_ab_1__23_), .ZN(u5_mult_82_n39) );
  AND2_X4 u5_mult_82_U131 ( .A1(u5_mult_82_ab_0__25_), .A2(
        u5_mult_82_ab_1__24_), .ZN(u5_mult_82_n38) );
  AND2_X4 u5_mult_82_U130 ( .A1(u5_mult_82_ab_0__26_), .A2(
        u5_mult_82_ab_1__25_), .ZN(u5_mult_82_n37) );
  AND2_X4 u5_mult_82_U129 ( .A1(u5_mult_82_ab_0__27_), .A2(
        u5_mult_82_ab_1__26_), .ZN(u5_mult_82_n36) );
  AND2_X4 u5_mult_82_U128 ( .A1(u5_mult_82_ab_0__28_), .A2(
        u5_mult_82_ab_1__27_), .ZN(u5_mult_82_n35) );
  AND2_X4 u5_mult_82_U127 ( .A1(u5_mult_82_ab_0__29_), .A2(
        u5_mult_82_ab_1__28_), .ZN(u5_mult_82_n34) );
  AND2_X4 u5_mult_82_U126 ( .A1(u5_mult_82_ab_0__4_), .A2(u5_mult_82_ab_1__3_), 
        .ZN(u5_mult_82_n33) );
  AND2_X4 u5_mult_82_U125 ( .A1(u5_mult_82_ab_0__5_), .A2(u5_mult_82_ab_1__4_), 
        .ZN(u5_mult_82_n32) );
  AND2_X4 u5_mult_82_U124 ( .A1(u5_mult_82_ab_0__7_), .A2(u5_mult_82_ab_1__6_), 
        .ZN(u5_mult_82_n31) );
  AND2_X4 u5_mult_82_U123 ( .A1(u5_mult_82_ab_0__9_), .A2(u5_mult_82_ab_1__8_), 
        .ZN(u5_mult_82_n30) );
  AND2_X4 u5_mult_82_U122 ( .A1(u5_mult_82_ab_0__2_), .A2(u5_mult_82_ab_1__1_), 
        .ZN(u5_mult_82_n29) );
  AND2_X4 u5_mult_82_U121 ( .A1(u5_mult_82_ab_0__3_), .A2(u5_mult_82_ab_1__2_), 
        .ZN(u5_mult_82_n28) );
  AND2_X4 u5_mult_82_U120 ( .A1(u5_mult_82_ab_0__30_), .A2(
        u5_mult_82_ab_1__29_), .ZN(u5_mult_82_n27) );
  AND2_X4 u5_mult_82_U119 ( .A1(u5_mult_82_ab_0__31_), .A2(
        u5_mult_82_ab_1__30_), .ZN(u5_mult_82_n26) );
  AND2_X4 u5_mult_82_U118 ( .A1(u5_mult_82_ab_0__32_), .A2(
        u5_mult_82_ab_1__31_), .ZN(u5_mult_82_n25) );
  AND2_X4 u5_mult_82_U117 ( .A1(u5_mult_82_ab_0__33_), .A2(
        u5_mult_82_ab_1__32_), .ZN(u5_mult_82_n24) );
  AND2_X4 u5_mult_82_U116 ( .A1(u5_mult_82_ab_0__34_), .A2(
        u5_mult_82_ab_1__33_), .ZN(u5_mult_82_n23) );
  AND2_X4 u5_mult_82_U115 ( .A1(u5_mult_82_ab_0__35_), .A2(
        u5_mult_82_ab_1__34_), .ZN(u5_mult_82_n22) );
  AND2_X4 u5_mult_82_U114 ( .A1(u5_mult_82_ab_0__36_), .A2(
        u5_mult_82_ab_1__35_), .ZN(u5_mult_82_n21) );
  AND2_X4 u5_mult_82_U113 ( .A1(u5_mult_82_ab_0__37_), .A2(
        u5_mult_82_ab_1__36_), .ZN(u5_mult_82_n20) );
  AND2_X4 u5_mult_82_U112 ( .A1(u5_mult_82_ab_0__38_), .A2(
        u5_mult_82_ab_1__37_), .ZN(u5_mult_82_n19) );
  AND2_X4 u5_mult_82_U111 ( .A1(u5_mult_82_ab_0__39_), .A2(
        u5_mult_82_ab_1__38_), .ZN(u5_mult_82_n18) );
  AND2_X4 u5_mult_82_U110 ( .A1(u5_mult_82_ab_0__40_), .A2(
        u5_mult_82_ab_1__39_), .ZN(u5_mult_82_n17) );
  AND2_X4 u5_mult_82_U109 ( .A1(u5_mult_82_ab_0__41_), .A2(
        u5_mult_82_ab_1__40_), .ZN(u5_mult_82_n16) );
  AND2_X4 u5_mult_82_U108 ( .A1(u5_mult_82_ab_0__42_), .A2(
        u5_mult_82_ab_1__41_), .ZN(u5_mult_82_n15) );
  AND2_X4 u5_mult_82_U107 ( .A1(u5_mult_82_ab_0__43_), .A2(
        u5_mult_82_ab_1__42_), .ZN(u5_mult_82_n14) );
  AND2_X4 u5_mult_82_U106 ( .A1(u5_mult_82_ab_0__44_), .A2(
        u5_mult_82_ab_1__43_), .ZN(u5_mult_82_n13) );
  AND2_X4 u5_mult_82_U105 ( .A1(u5_mult_82_ab_0__45_), .A2(
        u5_mult_82_ab_1__44_), .ZN(u5_mult_82_n12) );
  AND2_X4 u5_mult_82_U104 ( .A1(u5_mult_82_ab_0__46_), .A2(
        u5_mult_82_ab_1__45_), .ZN(u5_mult_82_n11) );
  AND2_X4 u5_mult_82_U103 ( .A1(u5_mult_82_ab_0__47_), .A2(
        u5_mult_82_ab_1__46_), .ZN(u5_mult_82_n10) );
  AND2_X4 u5_mult_82_U102 ( .A1(u5_mult_82_ab_0__48_), .A2(
        u5_mult_82_ab_1__47_), .ZN(u5_mult_82_n9) );
  AND2_X4 u5_mult_82_U101 ( .A1(u5_mult_82_ab_0__49_), .A2(
        u5_mult_82_ab_1__48_), .ZN(u5_mult_82_n8) );
  XOR2_X2 u5_mult_82_U100 ( .A(u5_mult_82_CARRYB_52__3_), .B(
        u5_mult_82_SUMB_52__4_), .Z(u5_mult_82_n7) );
  XOR2_X2 u5_mult_82_U99 ( .A(u5_mult_82_CARRYB_52__1_), .B(
        u5_mult_82_SUMB_52__2_), .Z(u5_mult_82_n6) );
  XOR2_X2 u5_mult_82_U98 ( .A(u5_mult_82_CARRYB_52__2_), .B(
        u5_mult_82_SUMB_52__3_), .Z(u5_mult_82_n5) );
  XOR2_X2 u5_mult_82_U97 ( .A(u5_mult_82_ab_1__51_), .B(u5_mult_82_ab_0__52_), 
        .Z(u5_mult_82_n4) );
  AND2_X4 u5_mult_82_U96 ( .A1(u5_mult_82_ab_0__50_), .A2(u5_mult_82_ab_1__49_), .ZN(u5_mult_82_n3) );
  INV_X4 u5_mult_82_U95 ( .A(fracta_mul[46]), .ZN(u5_mult_82_n224) );
  INV_X4 u5_mult_82_U94 ( .A(fracta_mul[50]), .ZN(u5_mult_82_n214) );
  INV_X4 u5_mult_82_U93 ( .A(n4602), .ZN(u5_mult_82_n449) );
  INV_X4 u5_mult_82_U92 ( .A(fracta_mul[41]), .ZN(u5_mult_82_n243) );
  INV_X4 u5_mult_82_U91 ( .A(fracta_mul[39]), .ZN(u5_mult_82_n248) );
  INV_X4 u5_mult_82_U90 ( .A(u5_mult_82_n454), .ZN(u5_mult_82_n235) );
  INV_X4 u5_mult_82_U89 ( .A(fracta_mul[35]), .ZN(u5_mult_82_n261) );
  INV_X4 u5_mult_82_U88 ( .A(fracta_mul[31]), .ZN(u5_mult_82_n269) );
  INV_X4 u5_mult_82_U87 ( .A(fracta_mul[28]), .ZN(u5_mult_82_n277) );
  INV_X4 u5_mult_82_U86 ( .A(fracta_mul[26]), .ZN(u5_mult_82_n281) );
  INV_X4 u5_mult_82_U85 ( .A(fracta_mul[18]), .ZN(u5_mult_82_n296) );
  INV_X4 u5_mult_82_U84 ( .A(u6_N2), .ZN(u5_mult_82_n442) );
  INV_X4 u5_mult_82_U83 ( .A(u6_N7), .ZN(u5_mult_82_n433) );
  INV_X4 u5_mult_82_U82 ( .A(u6_N9), .ZN(u5_mult_82_n429) );
  INV_X4 u5_mult_82_U81 ( .A(u6_N8), .ZN(u5_mult_82_n431) );
  INV_X4 u5_mult_82_U80 ( .A(fracta_mul[6]), .ZN(u5_mult_82_n316) );
  INV_X4 u5_mult_82_U79 ( .A(u6_N38), .ZN(u5_mult_82_n369) );
  INV_X4 u5_mult_82_U78 ( .A(u6_N11), .ZN(u5_mult_82_n426) );
  INV_X4 u5_mult_82_U77 ( .A(u6_N17), .ZN(u5_mult_82_n409) );
  INV_X4 u5_mult_82_U76 ( .A(u6_N32), .ZN(u5_mult_82_n379) );
  INV_X4 u5_mult_82_U75 ( .A(u6_N36), .ZN(u5_mult_82_n372) );
  INV_X4 u5_mult_82_U74 ( .A(u6_N19), .ZN(u5_mult_82_n404) );
  INV_X4 u5_mult_82_U73 ( .A(u6_N50), .ZN(u5_mult_82_n341) );
  INV_X4 u5_mult_82_U72 ( .A(u6_N52), .ZN(u5_mult_82_n337) );
  INV_X4 u5_mult_82_U71 ( .A(u6_N34), .ZN(u5_mult_82_n375) );
  INV_X4 u5_mult_82_U70 ( .A(u6_N43), .ZN(u5_mult_82_n356) );
  INV_X4 u5_mult_82_U69 ( .A(u6_N49), .ZN(u5_mult_82_n343) );
  INV_X4 u5_mult_82_U68 ( .A(u6_N51), .ZN(u5_mult_82_n339) );
  INV_X4 u5_mult_82_U67 ( .A(u6_N51), .ZN(u5_mult_82_n340) );
  INV_X4 u5_mult_82_U66 ( .A(fracta_mul[5]), .ZN(u5_mult_82_n319) );
  INV_X4 u5_mult_82_U65 ( .A(fracta_mul[1]), .ZN(u5_mult_82_n330) );
  INV_X4 u5_mult_82_U64 ( .A(fracta_mul[29]), .ZN(u5_mult_82_n274) );
  INV_X4 u5_mult_82_U63 ( .A(fracta_mul[21]), .ZN(u5_mult_82_n290) );
  INV_X4 u5_mult_82_U62 ( .A(fracta_mul[22]), .ZN(u5_mult_82_n288) );
  INV_X4 u5_mult_82_U61 ( .A(fracta_mul[24]), .ZN(u5_mult_82_n284) );
  INV_X4 u5_mult_82_U60 ( .A(fracta_mul[23]), .ZN(u5_mult_82_n286) );
  INV_X4 u5_mult_82_U59 ( .A(fracta_mul[20]), .ZN(u5_mult_82_n292) );
  INV_X4 u5_mult_82_U58 ( .A(fracta_mul[19]), .ZN(u5_mult_82_n293) );
  INV_X4 u5_mult_82_U57 ( .A(fracta_mul[7]), .ZN(u5_mult_82_n315) );
  INV_X4 u5_mult_82_U56 ( .A(u6_N5), .ZN(u5_mult_82_n437) );
  INV_X4 u5_mult_82_U55 ( .A(u6_N6), .ZN(u5_mult_82_n435) );
  INV_X4 u5_mult_82_U54 ( .A(u6_N4), .ZN(u5_mult_82_n439) );
  INV_X4 u5_mult_82_U53 ( .A(u6_N3), .ZN(u5_mult_82_n440) );
  INV_X4 u5_mult_82_U52 ( .A(u6_N10), .ZN(u5_mult_82_n427) );
  INV_X4 u5_mult_82_U51 ( .A(u6_N15), .ZN(u5_mult_82_n413) );
  INV_X4 u5_mult_82_U50 ( .A(u6_N16), .ZN(u5_mult_82_n410) );
  INV_X4 u5_mult_82_U49 ( .A(u6_N32), .ZN(u5_mult_82_n380) );
  INV_X4 u5_mult_82_U48 ( .A(u6_N37), .ZN(u5_mult_82_n370) );
  INV_X4 u5_mult_82_U47 ( .A(u6_N42), .ZN(u5_mult_82_n358) );
  INV_X4 u5_mult_82_U46 ( .A(u6_N44), .ZN(u5_mult_82_n353) );
  INV_X4 u5_mult_82_U45 ( .A(u6_N12), .ZN(u5_mult_82_n422) );
  INV_X4 u5_mult_82_U44 ( .A(u6_N14), .ZN(u5_mult_82_n416) );
  INV_X4 u5_mult_82_U43 ( .A(u6_N13), .ZN(u5_mult_82_n419) );
  INV_X4 u5_mult_82_U42 ( .A(u6_N35), .ZN(u5_mult_82_n373) );
  INV_X4 u5_mult_82_U41 ( .A(u6_N48), .ZN(u5_mult_82_n345) );
  INV_X4 u5_mult_82_U40 ( .A(u6_N47), .ZN(u5_mult_82_n347) );
  INV_X4 u5_mult_82_U39 ( .A(u6_N30), .ZN(u5_mult_82_n383) );
  INV_X4 u5_mult_82_U38 ( .A(u6_N41), .ZN(u5_mult_82_n361) );
  INV_X4 u5_mult_82_U37 ( .A(u6_N46), .ZN(u5_mult_82_n349) );
  INV_X4 u5_mult_82_U36 ( .A(u6_N31), .ZN(u5_mult_82_n381) );
  INV_X4 u5_mult_82_U35 ( .A(u6_N40), .ZN(u5_mult_82_n363) );
  INV_X4 u5_mult_82_U34 ( .A(u6_N45), .ZN(u5_mult_82_n351) );
  INV_X4 u5_mult_82_U33 ( .A(u6_N33), .ZN(u5_mult_82_n377) );
  INV_X4 u5_mult_82_U32 ( .A(u6_N39), .ZN(u5_mult_82_n365) );
  INV_X4 u5_mult_82_U31 ( .A(u6_N18), .ZN(u5_mult_82_n406) );
  INV_X4 u5_mult_82_U30 ( .A(u6_N51), .ZN(u5_mult_82_n338) );
  INV_X4 u5_mult_82_U29 ( .A(u6_N8), .ZN(u5_mult_82_n430) );
  INV_X4 u5_mult_82_U28 ( .A(fracta_mul[25]), .ZN(u5_mult_82_n282) );
  INV_X4 u5_mult_82_U27 ( .A(fracta_mul[14]), .ZN(u5_mult_82_n303) );
  INV_X4 u5_mult_82_U26 ( .A(u6_N0), .ZN(u5_mult_82_n446) );
  INV_X4 u5_mult_82_U25 ( .A(u6_N28), .ZN(u5_mult_82_n387) );
  INV_X4 u5_mult_82_U24 ( .A(u6_N5), .ZN(u5_mult_82_n436) );
  INV_X4 u5_mult_82_U23 ( .A(u6_N21), .ZN(u5_mult_82_n401) );
  INV_X4 u5_mult_82_U22 ( .A(u6_N22), .ZN(u5_mult_82_n399) );
  INV_X4 u5_mult_82_U21 ( .A(u6_N11), .ZN(u5_mult_82_n425) );
  INV_X4 u5_mult_82_U20 ( .A(u6_N17), .ZN(u5_mult_82_n408) );
  INV_X4 u5_mult_82_U19 ( .A(u6_N27), .ZN(u5_mult_82_n389) );
  INV_X4 u5_mult_82_U18 ( .A(u6_N24), .ZN(u5_mult_82_n395) );
  INV_X4 u5_mult_82_U17 ( .A(u6_N26), .ZN(u5_mult_82_n391) );
  INV_X4 u5_mult_82_U16 ( .A(u6_N7), .ZN(u5_mult_82_n432) );
  INV_X4 u5_mult_82_U15 ( .A(u6_N9), .ZN(u5_mult_82_n428) );
  INV_X4 u5_mult_82_U14 ( .A(u6_N4), .ZN(u5_mult_82_n438) );
  INV_X4 u5_mult_82_U13 ( .A(u6_N6), .ZN(u5_mult_82_n434) );
  INV_X4 u5_mult_82_U12 ( .A(fracta_mul[6]), .ZN(u5_mult_82_n317) );
  INV_X4 u5_mult_82_U11 ( .A(u6_N29), .ZN(u5_mult_82_n385) );
  INV_X4 u5_mult_82_U10 ( .A(u6_N23), .ZN(u5_mult_82_n397) );
  INV_X4 u5_mult_82_U9 ( .A(u6_N25), .ZN(u5_mult_82_n393) );
  INV_X4 u5_mult_82_U8 ( .A(u6_N52), .ZN(u5_mult_82_n336) );
  INV_X4 u5_mult_82_U7 ( .A(fracta_mul[16]), .ZN(u5_mult_82_n300) );
  INV_X4 u5_mult_82_U6 ( .A(fracta_mul[15]), .ZN(u5_mult_82_n302) );
  INV_X4 u5_mult_82_U5 ( .A(u6_N20), .ZN(u5_mult_82_n403) );
  INV_X4 u5_mult_82_U4 ( .A(fracta_mul[12]), .ZN(u5_mult_82_n307) );
  INV_X4 u5_mult_82_U3 ( .A(fracta_mul[13]), .ZN(u5_mult_82_n305) );
  INV_X4 u5_mult_82_U2 ( .A(fracta_mul[9]), .ZN(u5_mult_82_n311) );
  FA_X1 u5_mult_82_S3_2_51 ( .A(u5_mult_82_ab_2__51_), .B(u5_mult_82_n105), 
        .CI(u5_mult_82_ab_1__52_), .CO(u5_mult_82_CARRYB_2__51_), .S(
        u5_mult_82_SUMB_2__51_) );
  FA_X1 u5_mult_82_S2_2_50 ( .A(u5_mult_82_ab_2__50_), .B(u5_mult_82_n109), 
        .CI(u5_mult_82_n4), .CO(u5_mult_82_CARRYB_2__50_), .S(
        u5_mult_82_SUMB_2__50_) );
  FA_X1 u5_mult_82_S2_2_49 ( .A(u5_mult_82_ab_2__49_), .B(u5_mult_82_n3), .CI(
        u5_mult_82_n110), .CO(u5_mult_82_CARRYB_2__49_), .S(
        u5_mult_82_SUMB_2__49_) );
  FA_X1 u5_mult_82_S2_2_48 ( .A(u5_mult_82_ab_2__48_), .B(u5_mult_82_n8), .CI(
        u5_mult_82_n111), .CO(u5_mult_82_CARRYB_2__48_), .S(
        u5_mult_82_SUMB_2__48_) );
  FA_X1 u5_mult_82_S2_2_47 ( .A(u5_mult_82_ab_2__47_), .B(u5_mult_82_n9), .CI(
        u5_mult_82_n112), .CO(u5_mult_82_CARRYB_2__47_), .S(
        u5_mult_82_SUMB_2__47_) );
  FA_X1 u5_mult_82_S2_2_46 ( .A(u5_mult_82_ab_2__46_), .B(u5_mult_82_n10), 
        .CI(u5_mult_82_n113), .CO(u5_mult_82_CARRYB_2__46_), .S(
        u5_mult_82_SUMB_2__46_) );
  FA_X1 u5_mult_82_S2_2_45 ( .A(u5_mult_82_ab_2__45_), .B(u5_mult_82_n11), 
        .CI(u5_mult_82_n114), .CO(u5_mult_82_CARRYB_2__45_), .S(
        u5_mult_82_SUMB_2__45_) );
  FA_X1 u5_mult_82_S2_2_44 ( .A(u5_mult_82_ab_2__44_), .B(u5_mult_82_n12), 
        .CI(u5_mult_82_n115), .CO(u5_mult_82_CARRYB_2__44_), .S(
        u5_mult_82_SUMB_2__44_) );
  FA_X1 u5_mult_82_S2_2_43 ( .A(u5_mult_82_ab_2__43_), .B(u5_mult_82_n13), 
        .CI(u5_mult_82_n116), .CO(u5_mult_82_CARRYB_2__43_), .S(
        u5_mult_82_SUMB_2__43_) );
  FA_X1 u5_mult_82_S2_2_42 ( .A(u5_mult_82_ab_2__42_), .B(u5_mult_82_n14), 
        .CI(u5_mult_82_n117), .CO(u5_mult_82_CARRYB_2__42_), .S(
        u5_mult_82_SUMB_2__42_) );
  FA_X1 u5_mult_82_S2_2_41 ( .A(u5_mult_82_ab_2__41_), .B(u5_mult_82_n15), 
        .CI(u5_mult_82_n118), .CO(u5_mult_82_CARRYB_2__41_), .S(
        u5_mult_82_SUMB_2__41_) );
  FA_X1 u5_mult_82_S2_2_40 ( .A(u5_mult_82_ab_2__40_), .B(u5_mult_82_n16), 
        .CI(u5_mult_82_n119), .CO(u5_mult_82_CARRYB_2__40_), .S(
        u5_mult_82_SUMB_2__40_) );
  FA_X1 u5_mult_82_S2_2_39 ( .A(u5_mult_82_ab_2__39_), .B(u5_mult_82_n17), 
        .CI(u5_mult_82_n120), .CO(u5_mult_82_CARRYB_2__39_), .S(
        u5_mult_82_SUMB_2__39_) );
  FA_X1 u5_mult_82_S2_2_38 ( .A(u5_mult_82_ab_2__38_), .B(u5_mult_82_n18), 
        .CI(u5_mult_82_n121), .CO(u5_mult_82_CARRYB_2__38_), .S(
        u5_mult_82_SUMB_2__38_) );
  FA_X1 u5_mult_82_S2_2_37 ( .A(u5_mult_82_ab_2__37_), .B(u5_mult_82_n19), 
        .CI(u5_mult_82_n122), .CO(u5_mult_82_CARRYB_2__37_), .S(
        u5_mult_82_SUMB_2__37_) );
  FA_X1 u5_mult_82_S2_2_36 ( .A(u5_mult_82_ab_2__36_), .B(u5_mult_82_n20), 
        .CI(u5_mult_82_n123), .CO(u5_mult_82_CARRYB_2__36_), .S(
        u5_mult_82_SUMB_2__36_) );
  FA_X1 u5_mult_82_S2_2_35 ( .A(u5_mult_82_ab_2__35_), .B(u5_mult_82_n21), 
        .CI(u5_mult_82_n124), .CO(u5_mult_82_CARRYB_2__35_), .S(
        u5_mult_82_SUMB_2__35_) );
  FA_X1 u5_mult_82_S2_2_34 ( .A(u5_mult_82_ab_2__34_), .B(u5_mult_82_n22), 
        .CI(u5_mult_82_n125), .CO(u5_mult_82_CARRYB_2__34_), .S(
        u5_mult_82_SUMB_2__34_) );
  FA_X1 u5_mult_82_S2_2_33 ( .A(u5_mult_82_ab_2__33_), .B(u5_mult_82_n23), 
        .CI(u5_mult_82_n126), .CO(u5_mult_82_CARRYB_2__33_), .S(
        u5_mult_82_SUMB_2__33_) );
  FA_X1 u5_mult_82_S2_2_32 ( .A(u5_mult_82_ab_2__32_), .B(u5_mult_82_n24), 
        .CI(u5_mult_82_n127), .CO(u5_mult_82_CARRYB_2__32_), .S(
        u5_mult_82_SUMB_2__32_) );
  FA_X1 u5_mult_82_S2_2_31 ( .A(u5_mult_82_ab_2__31_), .B(u5_mult_82_n25), 
        .CI(u5_mult_82_n128), .CO(u5_mult_82_CARRYB_2__31_), .S(
        u5_mult_82_SUMB_2__31_) );
  FA_X1 u5_mult_82_S2_2_30 ( .A(u5_mult_82_ab_2__30_), .B(u5_mult_82_n26), 
        .CI(u5_mult_82_n129), .CO(u5_mult_82_CARRYB_2__30_), .S(
        u5_mult_82_SUMB_2__30_) );
  FA_X1 u5_mult_82_S2_2_29 ( .A(u5_mult_82_ab_2__29_), .B(u5_mult_82_n27), 
        .CI(u5_mult_82_n130), .CO(u5_mult_82_CARRYB_2__29_), .S(
        u5_mult_82_SUMB_2__29_) );
  FA_X1 u5_mult_82_S2_2_28 ( .A(u5_mult_82_ab_2__28_), .B(u5_mult_82_n34), 
        .CI(u5_mult_82_n131), .CO(u5_mult_82_CARRYB_2__28_), .S(
        u5_mult_82_SUMB_2__28_) );
  FA_X1 u5_mult_82_S2_2_27 ( .A(u5_mult_82_ab_2__27_), .B(u5_mult_82_n35), 
        .CI(u5_mult_82_n132), .CO(u5_mult_82_CARRYB_2__27_), .S(
        u5_mult_82_SUMB_2__27_) );
  FA_X1 u5_mult_82_S2_2_26 ( .A(u5_mult_82_ab_2__26_), .B(u5_mult_82_n36), 
        .CI(u5_mult_82_n133), .CO(u5_mult_82_CARRYB_2__26_), .S(
        u5_mult_82_SUMB_2__26_) );
  FA_X1 u5_mult_82_S2_2_25 ( .A(u5_mult_82_ab_2__25_), .B(u5_mult_82_n37), 
        .CI(u5_mult_82_n134), .CO(u5_mult_82_CARRYB_2__25_), .S(
        u5_mult_82_SUMB_2__25_) );
  FA_X1 u5_mult_82_S2_2_24 ( .A(u5_mult_82_ab_2__24_), .B(u5_mult_82_n38), 
        .CI(u5_mult_82_n135), .CO(u5_mult_82_CARRYB_2__24_), .S(
        u5_mult_82_SUMB_2__24_) );
  FA_X1 u5_mult_82_S2_2_23 ( .A(u5_mult_82_ab_2__23_), .B(u5_mult_82_n39), 
        .CI(u5_mult_82_n136), .CO(u5_mult_82_CARRYB_2__23_), .S(
        u5_mult_82_SUMB_2__23_) );
  FA_X1 u5_mult_82_S2_2_22 ( .A(u5_mult_82_ab_2__22_), .B(u5_mult_82_n40), 
        .CI(u5_mult_82_n137), .CO(u5_mult_82_CARRYB_2__22_), .S(
        u5_mult_82_SUMB_2__22_) );
  FA_X1 u5_mult_82_S2_2_21 ( .A(u5_mult_82_ab_2__21_), .B(u5_mult_82_n41), 
        .CI(u5_mult_82_n138), .CO(u5_mult_82_CARRYB_2__21_), .S(
        u5_mult_82_SUMB_2__21_) );
  FA_X1 u5_mult_82_S2_2_20 ( .A(u5_mult_82_ab_2__20_), .B(u5_mult_82_n42), 
        .CI(u5_mult_82_n139), .CO(u5_mult_82_CARRYB_2__20_), .S(
        u5_mult_82_SUMB_2__20_) );
  FA_X1 u5_mult_82_S2_2_19 ( .A(u5_mult_82_ab_2__19_), .B(u5_mult_82_n43), 
        .CI(u5_mult_82_n140), .CO(u5_mult_82_CARRYB_2__19_), .S(
        u5_mult_82_SUMB_2__19_) );
  FA_X1 u5_mult_82_S2_2_18 ( .A(u5_mult_82_ab_2__18_), .B(u5_mult_82_n44), 
        .CI(u5_mult_82_n141), .CO(u5_mult_82_CARRYB_2__18_), .S(
        u5_mult_82_SUMB_2__18_) );
  FA_X1 u5_mult_82_S2_2_17 ( .A(u5_mult_82_ab_2__17_), .B(u5_mult_82_n45), 
        .CI(u5_mult_82_n142), .CO(u5_mult_82_CARRYB_2__17_), .S(
        u5_mult_82_SUMB_2__17_) );
  FA_X1 u5_mult_82_S2_2_16 ( .A(u5_mult_82_ab_2__16_), .B(u5_mult_82_n46), 
        .CI(u5_mult_82_n143), .CO(u5_mult_82_CARRYB_2__16_), .S(
        u5_mult_82_SUMB_2__16_) );
  FA_X1 u5_mult_82_S2_2_15 ( .A(u5_mult_82_ab_2__15_), .B(u5_mult_82_n47), 
        .CI(u5_mult_82_n144), .CO(u5_mult_82_CARRYB_2__15_), .S(
        u5_mult_82_SUMB_2__15_) );
  FA_X1 u5_mult_82_S2_2_14 ( .A(u5_mult_82_ab_2__14_), .B(u5_mult_82_n48), 
        .CI(u5_mult_82_n145), .CO(u5_mult_82_CARRYB_2__14_), .S(
        u5_mult_82_SUMB_2__14_) );
  FA_X1 u5_mult_82_S2_2_13 ( .A(u5_mult_82_ab_2__13_), .B(u5_mult_82_n49), 
        .CI(u5_mult_82_n146), .CO(u5_mult_82_CARRYB_2__13_), .S(
        u5_mult_82_SUMB_2__13_) );
  FA_X1 u5_mult_82_S2_2_12 ( .A(u5_mult_82_ab_2__12_), .B(u5_mult_82_n50), 
        .CI(u5_mult_82_n147), .CO(u5_mult_82_CARRYB_2__12_), .S(
        u5_mult_82_SUMB_2__12_) );
  FA_X1 u5_mult_82_S2_2_11 ( .A(u5_mult_82_ab_2__11_), .B(u5_mult_82_n51), 
        .CI(u5_mult_82_n148), .CO(u5_mult_82_CARRYB_2__11_), .S(
        u5_mult_82_SUMB_2__11_) );
  FA_X1 u5_mult_82_S2_2_10 ( .A(u5_mult_82_ab_2__10_), .B(u5_mult_82_n52), 
        .CI(u5_mult_82_n149), .CO(u5_mult_82_CARRYB_2__10_), .S(
        u5_mult_82_SUMB_2__10_) );
  FA_X1 u5_mult_82_S2_2_9 ( .A(u5_mult_82_ab_2__9_), .B(u5_mult_82_n53), .CI(
        u5_mult_82_n150), .CO(u5_mult_82_CARRYB_2__9_), .S(
        u5_mult_82_SUMB_2__9_) );
  FA_X1 u5_mult_82_S2_2_8 ( .A(u5_mult_82_ab_2__8_), .B(u5_mult_82_n30), .CI(
        u5_mult_82_n151), .CO(u5_mult_82_CARRYB_2__8_), .S(
        u5_mult_82_SUMB_2__8_) );
  FA_X1 u5_mult_82_S2_2_7 ( .A(u5_mult_82_ab_2__7_), .B(u5_mult_82_n54), .CI(
        u5_mult_82_n152), .CO(u5_mult_82_CARRYB_2__7_), .S(
        u5_mult_82_SUMB_2__7_) );
  FA_X1 u5_mult_82_S2_2_6 ( .A(u5_mult_82_ab_2__6_), .B(u5_mult_82_n31), .CI(
        u5_mult_82_n153), .CO(u5_mult_82_CARRYB_2__6_), .S(
        u5_mult_82_SUMB_2__6_) );
  FA_X1 u5_mult_82_S2_2_5 ( .A(u5_mult_82_ab_2__5_), .B(u5_mult_82_n55), .CI(
        u5_mult_82_n154), .CO(u5_mult_82_CARRYB_2__5_), .S(
        u5_mult_82_SUMB_2__5_) );
  FA_X1 u5_mult_82_S2_2_4 ( .A(u5_mult_82_ab_2__4_), .B(u5_mult_82_n32), .CI(
        u5_mult_82_n155), .CO(u5_mult_82_CARRYB_2__4_), .S(
        u5_mult_82_SUMB_2__4_) );
  FA_X1 u5_mult_82_S2_2_3 ( .A(u5_mult_82_ab_2__3_), .B(u5_mult_82_n33), .CI(
        u5_mult_82_n156), .CO(u5_mult_82_CARRYB_2__3_), .S(
        u5_mult_82_SUMB_2__3_) );
  FA_X1 u5_mult_82_S2_2_2 ( .A(u5_mult_82_ab_2__2_), .B(u5_mult_82_n28), .CI(
        u5_mult_82_n157), .CO(u5_mult_82_CARRYB_2__2_), .S(
        u5_mult_82_SUMB_2__2_) );
  FA_X1 u5_mult_82_S2_2_1 ( .A(u5_mult_82_ab_2__1_), .B(u5_mult_82_n29), .CI(
        u5_mult_82_n158), .CO(u5_mult_82_CARRYB_2__1_), .S(
        u5_mult_82_SUMB_2__1_) );
  FA_X1 u5_mult_82_S1_2_0 ( .A(u5_mult_82_ab_2__0_), .B(u5_mult_82_n72), .CI(
        u5_mult_82_n171), .CO(u5_mult_82_CARRYB_2__0_), .S(u5_N2) );
  FA_X1 u5_mult_82_S3_3_51 ( .A(u5_mult_82_ab_3__51_), .B(
        u5_mult_82_CARRYB_2__51_), .CI(u5_mult_82_ab_2__52_), .CO(
        u5_mult_82_CARRYB_3__51_), .S(u5_mult_82_SUMB_3__51_) );
  FA_X1 u5_mult_82_S2_3_50 ( .A(u5_mult_82_ab_3__50_), .B(
        u5_mult_82_CARRYB_2__50_), .CI(u5_mult_82_SUMB_2__51_), .CO(
        u5_mult_82_CARRYB_3__50_), .S(u5_mult_82_SUMB_3__50_) );
  FA_X1 u5_mult_82_S2_3_49 ( .A(u5_mult_82_ab_3__49_), .B(
        u5_mult_82_CARRYB_2__49_), .CI(u5_mult_82_SUMB_2__50_), .CO(
        u5_mult_82_CARRYB_3__49_), .S(u5_mult_82_SUMB_3__49_) );
  FA_X1 u5_mult_82_S2_3_48 ( .A(u5_mult_82_ab_3__48_), .B(
        u5_mult_82_CARRYB_2__48_), .CI(u5_mult_82_SUMB_2__49_), .CO(
        u5_mult_82_CARRYB_3__48_), .S(u5_mult_82_SUMB_3__48_) );
  FA_X1 u5_mult_82_S2_3_47 ( .A(u5_mult_82_ab_3__47_), .B(
        u5_mult_82_CARRYB_2__47_), .CI(u5_mult_82_SUMB_2__48_), .CO(
        u5_mult_82_CARRYB_3__47_), .S(u5_mult_82_SUMB_3__47_) );
  FA_X1 u5_mult_82_S2_3_46 ( .A(u5_mult_82_ab_3__46_), .B(
        u5_mult_82_CARRYB_2__46_), .CI(u5_mult_82_SUMB_2__47_), .CO(
        u5_mult_82_CARRYB_3__46_), .S(u5_mult_82_SUMB_3__46_) );
  FA_X1 u5_mult_82_S2_3_45 ( .A(u5_mult_82_ab_3__45_), .B(
        u5_mult_82_CARRYB_2__45_), .CI(u5_mult_82_SUMB_2__46_), .CO(
        u5_mult_82_CARRYB_3__45_), .S(u5_mult_82_SUMB_3__45_) );
  FA_X1 u5_mult_82_S2_3_44 ( .A(u5_mult_82_ab_3__44_), .B(
        u5_mult_82_CARRYB_2__44_), .CI(u5_mult_82_SUMB_2__45_), .CO(
        u5_mult_82_CARRYB_3__44_), .S(u5_mult_82_SUMB_3__44_) );
  FA_X1 u5_mult_82_S2_3_43 ( .A(u5_mult_82_ab_3__43_), .B(
        u5_mult_82_CARRYB_2__43_), .CI(u5_mult_82_SUMB_2__44_), .CO(
        u5_mult_82_CARRYB_3__43_), .S(u5_mult_82_SUMB_3__43_) );
  FA_X1 u5_mult_82_S2_3_42 ( .A(u5_mult_82_ab_3__42_), .B(
        u5_mult_82_CARRYB_2__42_), .CI(u5_mult_82_SUMB_2__43_), .CO(
        u5_mult_82_CARRYB_3__42_), .S(u5_mult_82_SUMB_3__42_) );
  FA_X1 u5_mult_82_S2_3_41 ( .A(u5_mult_82_ab_3__41_), .B(
        u5_mult_82_CARRYB_2__41_), .CI(u5_mult_82_SUMB_2__42_), .CO(
        u5_mult_82_CARRYB_3__41_), .S(u5_mult_82_SUMB_3__41_) );
  FA_X1 u5_mult_82_S2_3_40 ( .A(u5_mult_82_ab_3__40_), .B(
        u5_mult_82_CARRYB_2__40_), .CI(u5_mult_82_SUMB_2__41_), .CO(
        u5_mult_82_CARRYB_3__40_), .S(u5_mult_82_SUMB_3__40_) );
  FA_X1 u5_mult_82_S2_3_39 ( .A(u5_mult_82_ab_3__39_), .B(
        u5_mult_82_CARRYB_2__39_), .CI(u5_mult_82_SUMB_2__40_), .CO(
        u5_mult_82_CARRYB_3__39_), .S(u5_mult_82_SUMB_3__39_) );
  FA_X1 u5_mult_82_S2_3_38 ( .A(u5_mult_82_ab_3__38_), .B(
        u5_mult_82_CARRYB_2__38_), .CI(u5_mult_82_SUMB_2__39_), .CO(
        u5_mult_82_CARRYB_3__38_), .S(u5_mult_82_SUMB_3__38_) );
  FA_X1 u5_mult_82_S2_3_37 ( .A(u5_mult_82_ab_3__37_), .B(
        u5_mult_82_CARRYB_2__37_), .CI(u5_mult_82_SUMB_2__38_), .CO(
        u5_mult_82_CARRYB_3__37_), .S(u5_mult_82_SUMB_3__37_) );
  FA_X1 u5_mult_82_S2_3_36 ( .A(u5_mult_82_ab_3__36_), .B(
        u5_mult_82_CARRYB_2__36_), .CI(u5_mult_82_SUMB_2__37_), .CO(
        u5_mult_82_CARRYB_3__36_), .S(u5_mult_82_SUMB_3__36_) );
  FA_X1 u5_mult_82_S2_3_35 ( .A(u5_mult_82_ab_3__35_), .B(
        u5_mult_82_CARRYB_2__35_), .CI(u5_mult_82_SUMB_2__36_), .CO(
        u5_mult_82_CARRYB_3__35_), .S(u5_mult_82_SUMB_3__35_) );
  FA_X1 u5_mult_82_S2_3_34 ( .A(u5_mult_82_ab_3__34_), .B(
        u5_mult_82_CARRYB_2__34_), .CI(u5_mult_82_SUMB_2__35_), .CO(
        u5_mult_82_CARRYB_3__34_), .S(u5_mult_82_SUMB_3__34_) );
  FA_X1 u5_mult_82_S2_3_33 ( .A(u5_mult_82_ab_3__33_), .B(
        u5_mult_82_CARRYB_2__33_), .CI(u5_mult_82_SUMB_2__34_), .CO(
        u5_mult_82_CARRYB_3__33_), .S(u5_mult_82_SUMB_3__33_) );
  FA_X1 u5_mult_82_S2_3_32 ( .A(u5_mult_82_ab_3__32_), .B(
        u5_mult_82_CARRYB_2__32_), .CI(u5_mult_82_SUMB_2__33_), .CO(
        u5_mult_82_CARRYB_3__32_), .S(u5_mult_82_SUMB_3__32_) );
  FA_X1 u5_mult_82_S2_3_31 ( .A(u5_mult_82_ab_3__31_), .B(
        u5_mult_82_CARRYB_2__31_), .CI(u5_mult_82_SUMB_2__32_), .CO(
        u5_mult_82_CARRYB_3__31_), .S(u5_mult_82_SUMB_3__31_) );
  FA_X1 u5_mult_82_S2_3_30 ( .A(u5_mult_82_ab_3__30_), .B(
        u5_mult_82_CARRYB_2__30_), .CI(u5_mult_82_SUMB_2__31_), .CO(
        u5_mult_82_CARRYB_3__30_), .S(u5_mult_82_SUMB_3__30_) );
  FA_X1 u5_mult_82_S2_3_29 ( .A(u5_mult_82_ab_3__29_), .B(
        u5_mult_82_CARRYB_2__29_), .CI(u5_mult_82_SUMB_2__30_), .CO(
        u5_mult_82_CARRYB_3__29_), .S(u5_mult_82_SUMB_3__29_) );
  FA_X1 u5_mult_82_S2_3_28 ( .A(u5_mult_82_ab_3__28_), .B(
        u5_mult_82_CARRYB_2__28_), .CI(u5_mult_82_SUMB_2__29_), .CO(
        u5_mult_82_CARRYB_3__28_), .S(u5_mult_82_SUMB_3__28_) );
  FA_X1 u5_mult_82_S2_3_27 ( .A(u5_mult_82_ab_3__27_), .B(
        u5_mult_82_CARRYB_2__27_), .CI(u5_mult_82_SUMB_2__28_), .CO(
        u5_mult_82_CARRYB_3__27_), .S(u5_mult_82_SUMB_3__27_) );
  FA_X1 u5_mult_82_S2_3_26 ( .A(u5_mult_82_ab_3__26_), .B(
        u5_mult_82_CARRYB_2__26_), .CI(u5_mult_82_SUMB_2__27_), .CO(
        u5_mult_82_CARRYB_3__26_), .S(u5_mult_82_SUMB_3__26_) );
  FA_X1 u5_mult_82_S2_3_25 ( .A(u5_mult_82_ab_3__25_), .B(
        u5_mult_82_CARRYB_2__25_), .CI(u5_mult_82_SUMB_2__26_), .CO(
        u5_mult_82_CARRYB_3__25_), .S(u5_mult_82_SUMB_3__25_) );
  FA_X1 u5_mult_82_S2_3_24 ( .A(u5_mult_82_ab_3__24_), .B(
        u5_mult_82_CARRYB_2__24_), .CI(u5_mult_82_SUMB_2__25_), .CO(
        u5_mult_82_CARRYB_3__24_), .S(u5_mult_82_SUMB_3__24_) );
  FA_X1 u5_mult_82_S2_3_23 ( .A(u5_mult_82_ab_3__23_), .B(
        u5_mult_82_CARRYB_2__23_), .CI(u5_mult_82_SUMB_2__24_), .CO(
        u5_mult_82_CARRYB_3__23_), .S(u5_mult_82_SUMB_3__23_) );
  FA_X1 u5_mult_82_S2_3_22 ( .A(u5_mult_82_ab_3__22_), .B(
        u5_mult_82_CARRYB_2__22_), .CI(u5_mult_82_SUMB_2__23_), .CO(
        u5_mult_82_CARRYB_3__22_), .S(u5_mult_82_SUMB_3__22_) );
  FA_X1 u5_mult_82_S2_3_21 ( .A(u5_mult_82_ab_3__21_), .B(
        u5_mult_82_CARRYB_2__21_), .CI(u5_mult_82_SUMB_2__22_), .CO(
        u5_mult_82_CARRYB_3__21_), .S(u5_mult_82_SUMB_3__21_) );
  FA_X1 u5_mult_82_S2_3_20 ( .A(u5_mult_82_ab_3__20_), .B(
        u5_mult_82_CARRYB_2__20_), .CI(u5_mult_82_SUMB_2__21_), .CO(
        u5_mult_82_CARRYB_3__20_), .S(u5_mult_82_SUMB_3__20_) );
  FA_X1 u5_mult_82_S2_3_19 ( .A(u5_mult_82_ab_3__19_), .B(
        u5_mult_82_CARRYB_2__19_), .CI(u5_mult_82_SUMB_2__20_), .CO(
        u5_mult_82_CARRYB_3__19_), .S(u5_mult_82_SUMB_3__19_) );
  FA_X1 u5_mult_82_S2_3_18 ( .A(u5_mult_82_ab_3__18_), .B(
        u5_mult_82_CARRYB_2__18_), .CI(u5_mult_82_SUMB_2__19_), .CO(
        u5_mult_82_CARRYB_3__18_), .S(u5_mult_82_SUMB_3__18_) );
  FA_X1 u5_mult_82_S2_3_17 ( .A(u5_mult_82_ab_3__17_), .B(
        u5_mult_82_CARRYB_2__17_), .CI(u5_mult_82_SUMB_2__18_), .CO(
        u5_mult_82_CARRYB_3__17_), .S(u5_mult_82_SUMB_3__17_) );
  FA_X1 u5_mult_82_S2_3_16 ( .A(u5_mult_82_ab_3__16_), .B(
        u5_mult_82_CARRYB_2__16_), .CI(u5_mult_82_SUMB_2__17_), .CO(
        u5_mult_82_CARRYB_3__16_), .S(u5_mult_82_SUMB_3__16_) );
  FA_X1 u5_mult_82_S2_3_15 ( .A(u5_mult_82_ab_3__15_), .B(
        u5_mult_82_CARRYB_2__15_), .CI(u5_mult_82_SUMB_2__16_), .CO(
        u5_mult_82_CARRYB_3__15_), .S(u5_mult_82_SUMB_3__15_) );
  FA_X1 u5_mult_82_S2_3_14 ( .A(u5_mult_82_ab_3__14_), .B(
        u5_mult_82_CARRYB_2__14_), .CI(u5_mult_82_SUMB_2__15_), .CO(
        u5_mult_82_CARRYB_3__14_), .S(u5_mult_82_SUMB_3__14_) );
  FA_X1 u5_mult_82_S2_3_13 ( .A(u5_mult_82_ab_3__13_), .B(
        u5_mult_82_CARRYB_2__13_), .CI(u5_mult_82_SUMB_2__14_), .CO(
        u5_mult_82_CARRYB_3__13_), .S(u5_mult_82_SUMB_3__13_) );
  FA_X1 u5_mult_82_S2_3_12 ( .A(u5_mult_82_ab_3__12_), .B(
        u5_mult_82_CARRYB_2__12_), .CI(u5_mult_82_SUMB_2__13_), .CO(
        u5_mult_82_CARRYB_3__12_), .S(u5_mult_82_SUMB_3__12_) );
  FA_X1 u5_mult_82_S2_3_11 ( .A(u5_mult_82_ab_3__11_), .B(
        u5_mult_82_CARRYB_2__11_), .CI(u5_mult_82_SUMB_2__12_), .CO(
        u5_mult_82_CARRYB_3__11_), .S(u5_mult_82_SUMB_3__11_) );
  FA_X1 u5_mult_82_S2_3_10 ( .A(u5_mult_82_ab_3__10_), .B(
        u5_mult_82_CARRYB_2__10_), .CI(u5_mult_82_SUMB_2__11_), .CO(
        u5_mult_82_CARRYB_3__10_), .S(u5_mult_82_SUMB_3__10_) );
  FA_X1 u5_mult_82_S2_3_9 ( .A(u5_mult_82_ab_3__9_), .B(
        u5_mult_82_CARRYB_2__9_), .CI(u5_mult_82_SUMB_2__10_), .CO(
        u5_mult_82_CARRYB_3__9_), .S(u5_mult_82_SUMB_3__9_) );
  FA_X1 u5_mult_82_S2_3_8 ( .A(u5_mult_82_ab_3__8_), .B(
        u5_mult_82_CARRYB_2__8_), .CI(u5_mult_82_SUMB_2__9_), .CO(
        u5_mult_82_CARRYB_3__8_), .S(u5_mult_82_SUMB_3__8_) );
  FA_X1 u5_mult_82_S2_3_7 ( .A(u5_mult_82_ab_3__7_), .B(
        u5_mult_82_CARRYB_2__7_), .CI(u5_mult_82_SUMB_2__8_), .CO(
        u5_mult_82_CARRYB_3__7_), .S(u5_mult_82_SUMB_3__7_) );
  FA_X1 u5_mult_82_S2_3_6 ( .A(u5_mult_82_ab_3__6_), .B(
        u5_mult_82_CARRYB_2__6_), .CI(u5_mult_82_SUMB_2__7_), .CO(
        u5_mult_82_CARRYB_3__6_), .S(u5_mult_82_SUMB_3__6_) );
  FA_X1 u5_mult_82_S2_3_5 ( .A(u5_mult_82_ab_3__5_), .B(
        u5_mult_82_CARRYB_2__5_), .CI(u5_mult_82_SUMB_2__6_), .CO(
        u5_mult_82_CARRYB_3__5_), .S(u5_mult_82_SUMB_3__5_) );
  FA_X1 u5_mult_82_S2_3_4 ( .A(u5_mult_82_ab_3__4_), .B(
        u5_mult_82_CARRYB_2__4_), .CI(u5_mult_82_SUMB_2__5_), .CO(
        u5_mult_82_CARRYB_3__4_), .S(u5_mult_82_SUMB_3__4_) );
  FA_X1 u5_mult_82_S2_3_3 ( .A(u5_mult_82_ab_3__3_), .B(
        u5_mult_82_CARRYB_2__3_), .CI(u5_mult_82_SUMB_2__4_), .CO(
        u5_mult_82_CARRYB_3__3_), .S(u5_mult_82_SUMB_3__3_) );
  FA_X1 u5_mult_82_S2_3_2 ( .A(u5_mult_82_ab_3__2_), .B(
        u5_mult_82_CARRYB_2__2_), .CI(u5_mult_82_SUMB_2__3_), .CO(
        u5_mult_82_CARRYB_3__2_), .S(u5_mult_82_SUMB_3__2_) );
  FA_X1 u5_mult_82_S2_3_1 ( .A(u5_mult_82_ab_3__1_), .B(
        u5_mult_82_CARRYB_2__1_), .CI(u5_mult_82_SUMB_2__2_), .CO(
        u5_mult_82_CARRYB_3__1_), .S(u5_mult_82_SUMB_3__1_) );
  FA_X1 u5_mult_82_S1_3_0 ( .A(u5_mult_82_ab_3__0_), .B(
        u5_mult_82_CARRYB_2__0_), .CI(u5_mult_82_SUMB_2__1_), .CO(
        u5_mult_82_CARRYB_3__0_), .S(u5_N3) );
  FA_X1 u5_mult_82_S3_4_51 ( .A(u5_mult_82_ab_4__51_), .B(
        u5_mult_82_CARRYB_3__51_), .CI(u5_mult_82_ab_3__52_), .CO(
        u5_mult_82_CARRYB_4__51_), .S(u5_mult_82_SUMB_4__51_) );
  FA_X1 u5_mult_82_S2_4_50 ( .A(u5_mult_82_ab_4__50_), .B(
        u5_mult_82_CARRYB_3__50_), .CI(u5_mult_82_SUMB_3__51_), .CO(
        u5_mult_82_CARRYB_4__50_), .S(u5_mult_82_SUMB_4__50_) );
  FA_X1 u5_mult_82_S2_4_49 ( .A(u5_mult_82_ab_4__49_), .B(
        u5_mult_82_CARRYB_3__49_), .CI(u5_mult_82_SUMB_3__50_), .CO(
        u5_mult_82_CARRYB_4__49_), .S(u5_mult_82_SUMB_4__49_) );
  FA_X1 u5_mult_82_S2_4_48 ( .A(u5_mult_82_ab_4__48_), .B(
        u5_mult_82_CARRYB_3__48_), .CI(u5_mult_82_SUMB_3__49_), .CO(
        u5_mult_82_CARRYB_4__48_), .S(u5_mult_82_SUMB_4__48_) );
  FA_X1 u5_mult_82_S2_4_47 ( .A(u5_mult_82_ab_4__47_), .B(
        u5_mult_82_CARRYB_3__47_), .CI(u5_mult_82_SUMB_3__48_), .CO(
        u5_mult_82_CARRYB_4__47_), .S(u5_mult_82_SUMB_4__47_) );
  FA_X1 u5_mult_82_S2_4_46 ( .A(u5_mult_82_ab_4__46_), .B(
        u5_mult_82_CARRYB_3__46_), .CI(u5_mult_82_SUMB_3__47_), .CO(
        u5_mult_82_CARRYB_4__46_), .S(u5_mult_82_SUMB_4__46_) );
  FA_X1 u5_mult_82_S2_4_45 ( .A(u5_mult_82_ab_4__45_), .B(
        u5_mult_82_CARRYB_3__45_), .CI(u5_mult_82_SUMB_3__46_), .CO(
        u5_mult_82_CARRYB_4__45_), .S(u5_mult_82_SUMB_4__45_) );
  FA_X1 u5_mult_82_S2_4_44 ( .A(u5_mult_82_ab_4__44_), .B(
        u5_mult_82_CARRYB_3__44_), .CI(u5_mult_82_SUMB_3__45_), .CO(
        u5_mult_82_CARRYB_4__44_), .S(u5_mult_82_SUMB_4__44_) );
  FA_X1 u5_mult_82_S2_4_43 ( .A(u5_mult_82_ab_4__43_), .B(
        u5_mult_82_CARRYB_3__43_), .CI(u5_mult_82_SUMB_3__44_), .CO(
        u5_mult_82_CARRYB_4__43_), .S(u5_mult_82_SUMB_4__43_) );
  FA_X1 u5_mult_82_S2_4_42 ( .A(u5_mult_82_ab_4__42_), .B(
        u5_mult_82_CARRYB_3__42_), .CI(u5_mult_82_SUMB_3__43_), .CO(
        u5_mult_82_CARRYB_4__42_), .S(u5_mult_82_SUMB_4__42_) );
  FA_X1 u5_mult_82_S2_4_41 ( .A(u5_mult_82_ab_4__41_), .B(
        u5_mult_82_CARRYB_3__41_), .CI(u5_mult_82_SUMB_3__42_), .CO(
        u5_mult_82_CARRYB_4__41_), .S(u5_mult_82_SUMB_4__41_) );
  FA_X1 u5_mult_82_S2_4_40 ( .A(u5_mult_82_ab_4__40_), .B(
        u5_mult_82_CARRYB_3__40_), .CI(u5_mult_82_SUMB_3__41_), .CO(
        u5_mult_82_CARRYB_4__40_), .S(u5_mult_82_SUMB_4__40_) );
  FA_X1 u5_mult_82_S2_4_39 ( .A(u5_mult_82_ab_4__39_), .B(
        u5_mult_82_CARRYB_3__39_), .CI(u5_mult_82_SUMB_3__40_), .CO(
        u5_mult_82_CARRYB_4__39_), .S(u5_mult_82_SUMB_4__39_) );
  FA_X1 u5_mult_82_S2_4_38 ( .A(u5_mult_82_ab_4__38_), .B(
        u5_mult_82_CARRYB_3__38_), .CI(u5_mult_82_SUMB_3__39_), .CO(
        u5_mult_82_CARRYB_4__38_), .S(u5_mult_82_SUMB_4__38_) );
  FA_X1 u5_mult_82_S2_4_37 ( .A(u5_mult_82_ab_4__37_), .B(
        u5_mult_82_CARRYB_3__37_), .CI(u5_mult_82_SUMB_3__38_), .CO(
        u5_mult_82_CARRYB_4__37_), .S(u5_mult_82_SUMB_4__37_) );
  FA_X1 u5_mult_82_S2_4_36 ( .A(u5_mult_82_ab_4__36_), .B(
        u5_mult_82_CARRYB_3__36_), .CI(u5_mult_82_SUMB_3__37_), .CO(
        u5_mult_82_CARRYB_4__36_), .S(u5_mult_82_SUMB_4__36_) );
  FA_X1 u5_mult_82_S2_4_35 ( .A(u5_mult_82_ab_4__35_), .B(
        u5_mult_82_CARRYB_3__35_), .CI(u5_mult_82_SUMB_3__36_), .CO(
        u5_mult_82_CARRYB_4__35_), .S(u5_mult_82_SUMB_4__35_) );
  FA_X1 u5_mult_82_S2_4_34 ( .A(u5_mult_82_ab_4__34_), .B(
        u5_mult_82_CARRYB_3__34_), .CI(u5_mult_82_SUMB_3__35_), .CO(
        u5_mult_82_CARRYB_4__34_), .S(u5_mult_82_SUMB_4__34_) );
  FA_X1 u5_mult_82_S2_4_33 ( .A(u5_mult_82_ab_4__33_), .B(
        u5_mult_82_CARRYB_3__33_), .CI(u5_mult_82_SUMB_3__34_), .CO(
        u5_mult_82_CARRYB_4__33_), .S(u5_mult_82_SUMB_4__33_) );
  FA_X1 u5_mult_82_S2_4_32 ( .A(u5_mult_82_ab_4__32_), .B(
        u5_mult_82_CARRYB_3__32_), .CI(u5_mult_82_SUMB_3__33_), .CO(
        u5_mult_82_CARRYB_4__32_), .S(u5_mult_82_SUMB_4__32_) );
  FA_X1 u5_mult_82_S2_4_31 ( .A(u5_mult_82_ab_4__31_), .B(
        u5_mult_82_CARRYB_3__31_), .CI(u5_mult_82_SUMB_3__32_), .CO(
        u5_mult_82_CARRYB_4__31_), .S(u5_mult_82_SUMB_4__31_) );
  FA_X1 u5_mult_82_S2_4_30 ( .A(u5_mult_82_ab_4__30_), .B(
        u5_mult_82_CARRYB_3__30_), .CI(u5_mult_82_SUMB_3__31_), .CO(
        u5_mult_82_CARRYB_4__30_), .S(u5_mult_82_SUMB_4__30_) );
  FA_X1 u5_mult_82_S2_4_29 ( .A(u5_mult_82_ab_4__29_), .B(
        u5_mult_82_CARRYB_3__29_), .CI(u5_mult_82_SUMB_3__30_), .CO(
        u5_mult_82_CARRYB_4__29_), .S(u5_mult_82_SUMB_4__29_) );
  FA_X1 u5_mult_82_S2_4_28 ( .A(u5_mult_82_ab_4__28_), .B(
        u5_mult_82_CARRYB_3__28_), .CI(u5_mult_82_SUMB_3__29_), .CO(
        u5_mult_82_CARRYB_4__28_), .S(u5_mult_82_SUMB_4__28_) );
  FA_X1 u5_mult_82_S2_4_27 ( .A(u5_mult_82_ab_4__27_), .B(
        u5_mult_82_CARRYB_3__27_), .CI(u5_mult_82_SUMB_3__28_), .CO(
        u5_mult_82_CARRYB_4__27_), .S(u5_mult_82_SUMB_4__27_) );
  FA_X1 u5_mult_82_S2_4_26 ( .A(u5_mult_82_ab_4__26_), .B(
        u5_mult_82_CARRYB_3__26_), .CI(u5_mult_82_SUMB_3__27_), .CO(
        u5_mult_82_CARRYB_4__26_), .S(u5_mult_82_SUMB_4__26_) );
  FA_X1 u5_mult_82_S2_4_25 ( .A(u5_mult_82_ab_4__25_), .B(
        u5_mult_82_CARRYB_3__25_), .CI(u5_mult_82_SUMB_3__26_), .CO(
        u5_mult_82_CARRYB_4__25_), .S(u5_mult_82_SUMB_4__25_) );
  FA_X1 u5_mult_82_S2_4_24 ( .A(u5_mult_82_ab_4__24_), .B(
        u5_mult_82_CARRYB_3__24_), .CI(u5_mult_82_SUMB_3__25_), .CO(
        u5_mult_82_CARRYB_4__24_), .S(u5_mult_82_SUMB_4__24_) );
  FA_X1 u5_mult_82_S2_4_23 ( .A(u5_mult_82_ab_4__23_), .B(
        u5_mult_82_CARRYB_3__23_), .CI(u5_mult_82_SUMB_3__24_), .CO(
        u5_mult_82_CARRYB_4__23_), .S(u5_mult_82_SUMB_4__23_) );
  FA_X1 u5_mult_82_S2_4_22 ( .A(u5_mult_82_ab_4__22_), .B(
        u5_mult_82_CARRYB_3__22_), .CI(u5_mult_82_SUMB_3__23_), .CO(
        u5_mult_82_CARRYB_4__22_), .S(u5_mult_82_SUMB_4__22_) );
  FA_X1 u5_mult_82_S2_4_21 ( .A(u5_mult_82_ab_4__21_), .B(
        u5_mult_82_CARRYB_3__21_), .CI(u5_mult_82_SUMB_3__22_), .CO(
        u5_mult_82_CARRYB_4__21_), .S(u5_mult_82_SUMB_4__21_) );
  FA_X1 u5_mult_82_S2_4_20 ( .A(u5_mult_82_ab_4__20_), .B(
        u5_mult_82_CARRYB_3__20_), .CI(u5_mult_82_SUMB_3__21_), .CO(
        u5_mult_82_CARRYB_4__20_), .S(u5_mult_82_SUMB_4__20_) );
  FA_X1 u5_mult_82_S2_4_19 ( .A(u5_mult_82_ab_4__19_), .B(
        u5_mult_82_CARRYB_3__19_), .CI(u5_mult_82_SUMB_3__20_), .CO(
        u5_mult_82_CARRYB_4__19_), .S(u5_mult_82_SUMB_4__19_) );
  FA_X1 u5_mult_82_S2_4_18 ( .A(u5_mult_82_ab_4__18_), .B(
        u5_mult_82_CARRYB_3__18_), .CI(u5_mult_82_SUMB_3__19_), .CO(
        u5_mult_82_CARRYB_4__18_), .S(u5_mult_82_SUMB_4__18_) );
  FA_X1 u5_mult_82_S2_4_17 ( .A(u5_mult_82_ab_4__17_), .B(
        u5_mult_82_CARRYB_3__17_), .CI(u5_mult_82_SUMB_3__18_), .CO(
        u5_mult_82_CARRYB_4__17_), .S(u5_mult_82_SUMB_4__17_) );
  FA_X1 u5_mult_82_S2_4_16 ( .A(u5_mult_82_ab_4__16_), .B(
        u5_mult_82_CARRYB_3__16_), .CI(u5_mult_82_SUMB_3__17_), .CO(
        u5_mult_82_CARRYB_4__16_), .S(u5_mult_82_SUMB_4__16_) );
  FA_X1 u5_mult_82_S2_4_15 ( .A(u5_mult_82_ab_4__15_), .B(
        u5_mult_82_CARRYB_3__15_), .CI(u5_mult_82_SUMB_3__16_), .CO(
        u5_mult_82_CARRYB_4__15_), .S(u5_mult_82_SUMB_4__15_) );
  FA_X1 u5_mult_82_S2_4_14 ( .A(u5_mult_82_ab_4__14_), .B(
        u5_mult_82_CARRYB_3__14_), .CI(u5_mult_82_SUMB_3__15_), .CO(
        u5_mult_82_CARRYB_4__14_), .S(u5_mult_82_SUMB_4__14_) );
  FA_X1 u5_mult_82_S2_4_13 ( .A(u5_mult_82_ab_4__13_), .B(
        u5_mult_82_CARRYB_3__13_), .CI(u5_mult_82_SUMB_3__14_), .CO(
        u5_mult_82_CARRYB_4__13_), .S(u5_mult_82_SUMB_4__13_) );
  FA_X1 u5_mult_82_S2_4_12 ( .A(u5_mult_82_ab_4__12_), .B(
        u5_mult_82_CARRYB_3__12_), .CI(u5_mult_82_SUMB_3__13_), .CO(
        u5_mult_82_CARRYB_4__12_), .S(u5_mult_82_SUMB_4__12_) );
  FA_X1 u5_mult_82_S2_4_11 ( .A(u5_mult_82_ab_4__11_), .B(
        u5_mult_82_CARRYB_3__11_), .CI(u5_mult_82_SUMB_3__12_), .CO(
        u5_mult_82_CARRYB_4__11_), .S(u5_mult_82_SUMB_4__11_) );
  FA_X1 u5_mult_82_S2_4_10 ( .A(u5_mult_82_ab_4__10_), .B(
        u5_mult_82_CARRYB_3__10_), .CI(u5_mult_82_SUMB_3__11_), .CO(
        u5_mult_82_CARRYB_4__10_), .S(u5_mult_82_SUMB_4__10_) );
  FA_X1 u5_mult_82_S2_4_9 ( .A(u5_mult_82_ab_4__9_), .B(
        u5_mult_82_CARRYB_3__9_), .CI(u5_mult_82_SUMB_3__10_), .CO(
        u5_mult_82_CARRYB_4__9_), .S(u5_mult_82_SUMB_4__9_) );
  FA_X1 u5_mult_82_S2_4_8 ( .A(u5_mult_82_ab_4__8_), .B(
        u5_mult_82_CARRYB_3__8_), .CI(u5_mult_82_SUMB_3__9_), .CO(
        u5_mult_82_CARRYB_4__8_), .S(u5_mult_82_SUMB_4__8_) );
  FA_X1 u5_mult_82_S2_4_7 ( .A(u5_mult_82_ab_4__7_), .B(
        u5_mult_82_CARRYB_3__7_), .CI(u5_mult_82_SUMB_3__8_), .CO(
        u5_mult_82_CARRYB_4__7_), .S(u5_mult_82_SUMB_4__7_) );
  FA_X1 u5_mult_82_S2_4_6 ( .A(u5_mult_82_ab_4__6_), .B(
        u5_mult_82_CARRYB_3__6_), .CI(u5_mult_82_SUMB_3__7_), .CO(
        u5_mult_82_CARRYB_4__6_), .S(u5_mult_82_SUMB_4__6_) );
  FA_X1 u5_mult_82_S2_4_5 ( .A(u5_mult_82_ab_4__5_), .B(
        u5_mult_82_CARRYB_3__5_), .CI(u5_mult_82_SUMB_3__6_), .CO(
        u5_mult_82_CARRYB_4__5_), .S(u5_mult_82_SUMB_4__5_) );
  FA_X1 u5_mult_82_S2_4_4 ( .A(u5_mult_82_ab_4__4_), .B(
        u5_mult_82_CARRYB_3__4_), .CI(u5_mult_82_SUMB_3__5_), .CO(
        u5_mult_82_CARRYB_4__4_), .S(u5_mult_82_SUMB_4__4_) );
  FA_X1 u5_mult_82_S2_4_3 ( .A(u5_mult_82_ab_4__3_), .B(
        u5_mult_82_CARRYB_3__3_), .CI(u5_mult_82_SUMB_3__4_), .CO(
        u5_mult_82_CARRYB_4__3_), .S(u5_mult_82_SUMB_4__3_) );
  FA_X1 u5_mult_82_S2_4_2 ( .A(u5_mult_82_ab_4__2_), .B(
        u5_mult_82_CARRYB_3__2_), .CI(u5_mult_82_SUMB_3__3_), .CO(
        u5_mult_82_CARRYB_4__2_), .S(u5_mult_82_SUMB_4__2_) );
  FA_X1 u5_mult_82_S2_4_1 ( .A(u5_mult_82_ab_4__1_), .B(
        u5_mult_82_CARRYB_3__1_), .CI(u5_mult_82_SUMB_3__2_), .CO(
        u5_mult_82_CARRYB_4__1_), .S(u5_mult_82_SUMB_4__1_) );
  FA_X1 u5_mult_82_S1_4_0 ( .A(u5_mult_82_ab_4__0_), .B(
        u5_mult_82_CARRYB_3__0_), .CI(u5_mult_82_SUMB_3__1_), .CO(
        u5_mult_82_CARRYB_4__0_), .S(u5_N4) );
  FA_X1 u5_mult_82_S3_5_51 ( .A(u5_mult_82_ab_5__51_), .B(
        u5_mult_82_CARRYB_4__51_), .CI(u5_mult_82_ab_4__52_), .CO(
        u5_mult_82_CARRYB_5__51_), .S(u5_mult_82_SUMB_5__51_) );
  FA_X1 u5_mult_82_S2_5_50 ( .A(u5_mult_82_ab_5__50_), .B(
        u5_mult_82_CARRYB_4__50_), .CI(u5_mult_82_SUMB_4__51_), .CO(
        u5_mult_82_CARRYB_5__50_), .S(u5_mult_82_SUMB_5__50_) );
  FA_X1 u5_mult_82_S2_5_49 ( .A(u5_mult_82_ab_5__49_), .B(
        u5_mult_82_CARRYB_4__49_), .CI(u5_mult_82_SUMB_4__50_), .CO(
        u5_mult_82_CARRYB_5__49_), .S(u5_mult_82_SUMB_5__49_) );
  FA_X1 u5_mult_82_S2_5_48 ( .A(u5_mult_82_ab_5__48_), .B(
        u5_mult_82_CARRYB_4__48_), .CI(u5_mult_82_SUMB_4__49_), .CO(
        u5_mult_82_CARRYB_5__48_), .S(u5_mult_82_SUMB_5__48_) );
  FA_X1 u5_mult_82_S2_5_47 ( .A(u5_mult_82_ab_5__47_), .B(
        u5_mult_82_CARRYB_4__47_), .CI(u5_mult_82_SUMB_4__48_), .CO(
        u5_mult_82_CARRYB_5__47_), .S(u5_mult_82_SUMB_5__47_) );
  FA_X1 u5_mult_82_S2_5_46 ( .A(u5_mult_82_ab_5__46_), .B(
        u5_mult_82_CARRYB_4__46_), .CI(u5_mult_82_SUMB_4__47_), .CO(
        u5_mult_82_CARRYB_5__46_), .S(u5_mult_82_SUMB_5__46_) );
  FA_X1 u5_mult_82_S2_5_45 ( .A(u5_mult_82_ab_5__45_), .B(
        u5_mult_82_CARRYB_4__45_), .CI(u5_mult_82_SUMB_4__46_), .CO(
        u5_mult_82_CARRYB_5__45_), .S(u5_mult_82_SUMB_5__45_) );
  FA_X1 u5_mult_82_S2_5_44 ( .A(u5_mult_82_ab_5__44_), .B(
        u5_mult_82_CARRYB_4__44_), .CI(u5_mult_82_SUMB_4__45_), .CO(
        u5_mult_82_CARRYB_5__44_), .S(u5_mult_82_SUMB_5__44_) );
  FA_X1 u5_mult_82_S2_5_43 ( .A(u5_mult_82_ab_5__43_), .B(
        u5_mult_82_CARRYB_4__43_), .CI(u5_mult_82_SUMB_4__44_), .CO(
        u5_mult_82_CARRYB_5__43_), .S(u5_mult_82_SUMB_5__43_) );
  FA_X1 u5_mult_82_S2_5_42 ( .A(u5_mult_82_ab_5__42_), .B(
        u5_mult_82_CARRYB_4__42_), .CI(u5_mult_82_SUMB_4__43_), .CO(
        u5_mult_82_CARRYB_5__42_), .S(u5_mult_82_SUMB_5__42_) );
  FA_X1 u5_mult_82_S2_5_41 ( .A(u5_mult_82_ab_5__41_), .B(
        u5_mult_82_CARRYB_4__41_), .CI(u5_mult_82_SUMB_4__42_), .CO(
        u5_mult_82_CARRYB_5__41_), .S(u5_mult_82_SUMB_5__41_) );
  FA_X1 u5_mult_82_S2_5_40 ( .A(u5_mult_82_ab_5__40_), .B(
        u5_mult_82_CARRYB_4__40_), .CI(u5_mult_82_SUMB_4__41_), .CO(
        u5_mult_82_CARRYB_5__40_), .S(u5_mult_82_SUMB_5__40_) );
  FA_X1 u5_mult_82_S2_5_39 ( .A(u5_mult_82_ab_5__39_), .B(
        u5_mult_82_CARRYB_4__39_), .CI(u5_mult_82_SUMB_4__40_), .CO(
        u5_mult_82_CARRYB_5__39_), .S(u5_mult_82_SUMB_5__39_) );
  FA_X1 u5_mult_82_S2_5_38 ( .A(u5_mult_82_ab_5__38_), .B(
        u5_mult_82_CARRYB_4__38_), .CI(u5_mult_82_SUMB_4__39_), .CO(
        u5_mult_82_CARRYB_5__38_), .S(u5_mult_82_SUMB_5__38_) );
  FA_X1 u5_mult_82_S2_5_37 ( .A(u5_mult_82_ab_5__37_), .B(
        u5_mult_82_CARRYB_4__37_), .CI(u5_mult_82_SUMB_4__38_), .CO(
        u5_mult_82_CARRYB_5__37_), .S(u5_mult_82_SUMB_5__37_) );
  FA_X1 u5_mult_82_S2_5_36 ( .A(u5_mult_82_ab_5__36_), .B(
        u5_mult_82_CARRYB_4__36_), .CI(u5_mult_82_SUMB_4__37_), .CO(
        u5_mult_82_CARRYB_5__36_), .S(u5_mult_82_SUMB_5__36_) );
  FA_X1 u5_mult_82_S2_5_35 ( .A(u5_mult_82_ab_5__35_), .B(
        u5_mult_82_CARRYB_4__35_), .CI(u5_mult_82_SUMB_4__36_), .CO(
        u5_mult_82_CARRYB_5__35_), .S(u5_mult_82_SUMB_5__35_) );
  FA_X1 u5_mult_82_S2_5_34 ( .A(u5_mult_82_ab_5__34_), .B(
        u5_mult_82_CARRYB_4__34_), .CI(u5_mult_82_SUMB_4__35_), .CO(
        u5_mult_82_CARRYB_5__34_), .S(u5_mult_82_SUMB_5__34_) );
  FA_X1 u5_mult_82_S2_5_33 ( .A(u5_mult_82_ab_5__33_), .B(
        u5_mult_82_CARRYB_4__33_), .CI(u5_mult_82_SUMB_4__34_), .CO(
        u5_mult_82_CARRYB_5__33_), .S(u5_mult_82_SUMB_5__33_) );
  FA_X1 u5_mult_82_S2_5_32 ( .A(u5_mult_82_ab_5__32_), .B(
        u5_mult_82_CARRYB_4__32_), .CI(u5_mult_82_SUMB_4__33_), .CO(
        u5_mult_82_CARRYB_5__32_), .S(u5_mult_82_SUMB_5__32_) );
  FA_X1 u5_mult_82_S2_5_31 ( .A(u5_mult_82_ab_5__31_), .B(
        u5_mult_82_CARRYB_4__31_), .CI(u5_mult_82_SUMB_4__32_), .CO(
        u5_mult_82_CARRYB_5__31_), .S(u5_mult_82_SUMB_5__31_) );
  FA_X1 u5_mult_82_S2_5_30 ( .A(u5_mult_82_ab_5__30_), .B(
        u5_mult_82_CARRYB_4__30_), .CI(u5_mult_82_SUMB_4__31_), .CO(
        u5_mult_82_CARRYB_5__30_), .S(u5_mult_82_SUMB_5__30_) );
  FA_X1 u5_mult_82_S2_5_29 ( .A(u5_mult_82_ab_5__29_), .B(
        u5_mult_82_CARRYB_4__29_), .CI(u5_mult_82_SUMB_4__30_), .CO(
        u5_mult_82_CARRYB_5__29_), .S(u5_mult_82_SUMB_5__29_) );
  FA_X1 u5_mult_82_S2_5_28 ( .A(u5_mult_82_ab_5__28_), .B(
        u5_mult_82_CARRYB_4__28_), .CI(u5_mult_82_SUMB_4__29_), .CO(
        u5_mult_82_CARRYB_5__28_), .S(u5_mult_82_SUMB_5__28_) );
  FA_X1 u5_mult_82_S2_5_27 ( .A(u5_mult_82_ab_5__27_), .B(
        u5_mult_82_CARRYB_4__27_), .CI(u5_mult_82_SUMB_4__28_), .CO(
        u5_mult_82_CARRYB_5__27_), .S(u5_mult_82_SUMB_5__27_) );
  FA_X1 u5_mult_82_S2_5_26 ( .A(u5_mult_82_ab_5__26_), .B(
        u5_mult_82_CARRYB_4__26_), .CI(u5_mult_82_SUMB_4__27_), .CO(
        u5_mult_82_CARRYB_5__26_), .S(u5_mult_82_SUMB_5__26_) );
  FA_X1 u5_mult_82_S2_5_25 ( .A(u5_mult_82_ab_5__25_), .B(
        u5_mult_82_CARRYB_4__25_), .CI(u5_mult_82_SUMB_4__26_), .CO(
        u5_mult_82_CARRYB_5__25_), .S(u5_mult_82_SUMB_5__25_) );
  FA_X1 u5_mult_82_S2_5_24 ( .A(u5_mult_82_ab_5__24_), .B(
        u5_mult_82_CARRYB_4__24_), .CI(u5_mult_82_SUMB_4__25_), .CO(
        u5_mult_82_CARRYB_5__24_), .S(u5_mult_82_SUMB_5__24_) );
  FA_X1 u5_mult_82_S2_5_23 ( .A(u5_mult_82_ab_5__23_), .B(
        u5_mult_82_CARRYB_4__23_), .CI(u5_mult_82_SUMB_4__24_), .CO(
        u5_mult_82_CARRYB_5__23_), .S(u5_mult_82_SUMB_5__23_) );
  FA_X1 u5_mult_82_S2_5_22 ( .A(u5_mult_82_ab_5__22_), .B(
        u5_mult_82_CARRYB_4__22_), .CI(u5_mult_82_SUMB_4__23_), .CO(
        u5_mult_82_CARRYB_5__22_), .S(u5_mult_82_SUMB_5__22_) );
  FA_X1 u5_mult_82_S2_5_21 ( .A(u5_mult_82_ab_5__21_), .B(
        u5_mult_82_CARRYB_4__21_), .CI(u5_mult_82_SUMB_4__22_), .CO(
        u5_mult_82_CARRYB_5__21_), .S(u5_mult_82_SUMB_5__21_) );
  FA_X1 u5_mult_82_S2_5_20 ( .A(u5_mult_82_ab_5__20_), .B(
        u5_mult_82_CARRYB_4__20_), .CI(u5_mult_82_SUMB_4__21_), .CO(
        u5_mult_82_CARRYB_5__20_), .S(u5_mult_82_SUMB_5__20_) );
  FA_X1 u5_mult_82_S2_5_19 ( .A(u5_mult_82_ab_5__19_), .B(
        u5_mult_82_CARRYB_4__19_), .CI(u5_mult_82_SUMB_4__20_), .CO(
        u5_mult_82_CARRYB_5__19_), .S(u5_mult_82_SUMB_5__19_) );
  FA_X1 u5_mult_82_S2_5_18 ( .A(u5_mult_82_ab_5__18_), .B(
        u5_mult_82_CARRYB_4__18_), .CI(u5_mult_82_SUMB_4__19_), .CO(
        u5_mult_82_CARRYB_5__18_), .S(u5_mult_82_SUMB_5__18_) );
  FA_X1 u5_mult_82_S2_5_17 ( .A(u5_mult_82_ab_5__17_), .B(
        u5_mult_82_CARRYB_4__17_), .CI(u5_mult_82_SUMB_4__18_), .CO(
        u5_mult_82_CARRYB_5__17_), .S(u5_mult_82_SUMB_5__17_) );
  FA_X1 u5_mult_82_S2_5_16 ( .A(u5_mult_82_ab_5__16_), .B(
        u5_mult_82_CARRYB_4__16_), .CI(u5_mult_82_SUMB_4__17_), .CO(
        u5_mult_82_CARRYB_5__16_), .S(u5_mult_82_SUMB_5__16_) );
  FA_X1 u5_mult_82_S2_5_15 ( .A(u5_mult_82_ab_5__15_), .B(
        u5_mult_82_CARRYB_4__15_), .CI(u5_mult_82_SUMB_4__16_), .CO(
        u5_mult_82_CARRYB_5__15_), .S(u5_mult_82_SUMB_5__15_) );
  FA_X1 u5_mult_82_S2_5_14 ( .A(u5_mult_82_ab_5__14_), .B(
        u5_mult_82_CARRYB_4__14_), .CI(u5_mult_82_SUMB_4__15_), .CO(
        u5_mult_82_CARRYB_5__14_), .S(u5_mult_82_SUMB_5__14_) );
  FA_X1 u5_mult_82_S2_5_13 ( .A(u5_mult_82_ab_5__13_), .B(
        u5_mult_82_CARRYB_4__13_), .CI(u5_mult_82_SUMB_4__14_), .CO(
        u5_mult_82_CARRYB_5__13_), .S(u5_mult_82_SUMB_5__13_) );
  FA_X1 u5_mult_82_S2_5_12 ( .A(u5_mult_82_ab_5__12_), .B(
        u5_mult_82_CARRYB_4__12_), .CI(u5_mult_82_SUMB_4__13_), .CO(
        u5_mult_82_CARRYB_5__12_), .S(u5_mult_82_SUMB_5__12_) );
  FA_X1 u5_mult_82_S2_5_11 ( .A(u5_mult_82_ab_5__11_), .B(
        u5_mult_82_CARRYB_4__11_), .CI(u5_mult_82_SUMB_4__12_), .CO(
        u5_mult_82_CARRYB_5__11_), .S(u5_mult_82_SUMB_5__11_) );
  FA_X1 u5_mult_82_S2_5_10 ( .A(u5_mult_82_ab_5__10_), .B(
        u5_mult_82_CARRYB_4__10_), .CI(u5_mult_82_SUMB_4__11_), .CO(
        u5_mult_82_CARRYB_5__10_), .S(u5_mult_82_SUMB_5__10_) );
  FA_X1 u5_mult_82_S2_5_9 ( .A(u5_mult_82_ab_5__9_), .B(
        u5_mult_82_CARRYB_4__9_), .CI(u5_mult_82_SUMB_4__10_), .CO(
        u5_mult_82_CARRYB_5__9_), .S(u5_mult_82_SUMB_5__9_) );
  FA_X1 u5_mult_82_S2_5_8 ( .A(u5_mult_82_ab_5__8_), .B(
        u5_mult_82_CARRYB_4__8_), .CI(u5_mult_82_SUMB_4__9_), .CO(
        u5_mult_82_CARRYB_5__8_), .S(u5_mult_82_SUMB_5__8_) );
  FA_X1 u5_mult_82_S2_5_7 ( .A(u5_mult_82_ab_5__7_), .B(
        u5_mult_82_CARRYB_4__7_), .CI(u5_mult_82_SUMB_4__8_), .CO(
        u5_mult_82_CARRYB_5__7_), .S(u5_mult_82_SUMB_5__7_) );
  FA_X1 u5_mult_82_S2_5_6 ( .A(u5_mult_82_ab_5__6_), .B(
        u5_mult_82_CARRYB_4__6_), .CI(u5_mult_82_SUMB_4__7_), .CO(
        u5_mult_82_CARRYB_5__6_), .S(u5_mult_82_SUMB_5__6_) );
  FA_X1 u5_mult_82_S2_5_5 ( .A(u5_mult_82_ab_5__5_), .B(
        u5_mult_82_CARRYB_4__5_), .CI(u5_mult_82_SUMB_4__6_), .CO(
        u5_mult_82_CARRYB_5__5_), .S(u5_mult_82_SUMB_5__5_) );
  FA_X1 u5_mult_82_S2_5_4 ( .A(u5_mult_82_ab_5__4_), .B(
        u5_mult_82_CARRYB_4__4_), .CI(u5_mult_82_SUMB_4__5_), .CO(
        u5_mult_82_CARRYB_5__4_), .S(u5_mult_82_SUMB_5__4_) );
  FA_X1 u5_mult_82_S2_5_3 ( .A(u5_mult_82_ab_5__3_), .B(
        u5_mult_82_CARRYB_4__3_), .CI(u5_mult_82_SUMB_4__4_), .CO(
        u5_mult_82_CARRYB_5__3_), .S(u5_mult_82_SUMB_5__3_) );
  FA_X1 u5_mult_82_S2_5_2 ( .A(u5_mult_82_ab_5__2_), .B(
        u5_mult_82_CARRYB_4__2_), .CI(u5_mult_82_SUMB_4__3_), .CO(
        u5_mult_82_CARRYB_5__2_), .S(u5_mult_82_SUMB_5__2_) );
  FA_X1 u5_mult_82_S2_5_1 ( .A(u5_mult_82_ab_5__1_), .B(
        u5_mult_82_CARRYB_4__1_), .CI(u5_mult_82_SUMB_4__2_), .CO(
        u5_mult_82_CARRYB_5__1_), .S(u5_mult_82_SUMB_5__1_) );
  FA_X1 u5_mult_82_S1_5_0 ( .A(u5_mult_82_ab_5__0_), .B(
        u5_mult_82_CARRYB_4__0_), .CI(u5_mult_82_SUMB_4__1_), .CO(
        u5_mult_82_CARRYB_5__0_), .S(u5_N5) );
  FA_X1 u5_mult_82_S3_6_51 ( .A(u5_mult_82_ab_6__51_), .B(
        u5_mult_82_CARRYB_5__51_), .CI(u5_mult_82_ab_5__52_), .CO(
        u5_mult_82_CARRYB_6__51_), .S(u5_mult_82_SUMB_6__51_) );
  FA_X1 u5_mult_82_S2_6_50 ( .A(u5_mult_82_ab_6__50_), .B(
        u5_mult_82_CARRYB_5__50_), .CI(u5_mult_82_SUMB_5__51_), .CO(
        u5_mult_82_CARRYB_6__50_), .S(u5_mult_82_SUMB_6__50_) );
  FA_X1 u5_mult_82_S2_6_49 ( .A(u5_mult_82_ab_6__49_), .B(
        u5_mult_82_CARRYB_5__49_), .CI(u5_mult_82_SUMB_5__50_), .CO(
        u5_mult_82_CARRYB_6__49_), .S(u5_mult_82_SUMB_6__49_) );
  FA_X1 u5_mult_82_S2_6_48 ( .A(u5_mult_82_ab_6__48_), .B(
        u5_mult_82_CARRYB_5__48_), .CI(u5_mult_82_SUMB_5__49_), .CO(
        u5_mult_82_CARRYB_6__48_), .S(u5_mult_82_SUMB_6__48_) );
  FA_X1 u5_mult_82_S2_6_47 ( .A(u5_mult_82_ab_6__47_), .B(
        u5_mult_82_CARRYB_5__47_), .CI(u5_mult_82_SUMB_5__48_), .CO(
        u5_mult_82_CARRYB_6__47_), .S(u5_mult_82_SUMB_6__47_) );
  FA_X1 u5_mult_82_S2_6_46 ( .A(u5_mult_82_ab_6__46_), .B(
        u5_mult_82_CARRYB_5__46_), .CI(u5_mult_82_SUMB_5__47_), .CO(
        u5_mult_82_CARRYB_6__46_), .S(u5_mult_82_SUMB_6__46_) );
  FA_X1 u5_mult_82_S2_6_45 ( .A(u5_mult_82_ab_6__45_), .B(
        u5_mult_82_CARRYB_5__45_), .CI(u5_mult_82_SUMB_5__46_), .CO(
        u5_mult_82_CARRYB_6__45_), .S(u5_mult_82_SUMB_6__45_) );
  FA_X1 u5_mult_82_S2_6_44 ( .A(u5_mult_82_ab_6__44_), .B(
        u5_mult_82_CARRYB_5__44_), .CI(u5_mult_82_SUMB_5__45_), .CO(
        u5_mult_82_CARRYB_6__44_), .S(u5_mult_82_SUMB_6__44_) );
  FA_X1 u5_mult_82_S2_6_43 ( .A(u5_mult_82_ab_6__43_), .B(
        u5_mult_82_CARRYB_5__43_), .CI(u5_mult_82_SUMB_5__44_), .CO(
        u5_mult_82_CARRYB_6__43_), .S(u5_mult_82_SUMB_6__43_) );
  FA_X1 u5_mult_82_S2_6_42 ( .A(u5_mult_82_ab_6__42_), .B(
        u5_mult_82_CARRYB_5__42_), .CI(u5_mult_82_SUMB_5__43_), .CO(
        u5_mult_82_CARRYB_6__42_), .S(u5_mult_82_SUMB_6__42_) );
  FA_X1 u5_mult_82_S2_6_41 ( .A(u5_mult_82_ab_6__41_), .B(
        u5_mult_82_CARRYB_5__41_), .CI(u5_mult_82_SUMB_5__42_), .CO(
        u5_mult_82_CARRYB_6__41_), .S(u5_mult_82_SUMB_6__41_) );
  FA_X1 u5_mult_82_S2_6_40 ( .A(u5_mult_82_ab_6__40_), .B(
        u5_mult_82_CARRYB_5__40_), .CI(u5_mult_82_SUMB_5__41_), .CO(
        u5_mult_82_CARRYB_6__40_), .S(u5_mult_82_SUMB_6__40_) );
  FA_X1 u5_mult_82_S2_6_39 ( .A(u5_mult_82_ab_6__39_), .B(
        u5_mult_82_CARRYB_5__39_), .CI(u5_mult_82_SUMB_5__40_), .CO(
        u5_mult_82_CARRYB_6__39_), .S(u5_mult_82_SUMB_6__39_) );
  FA_X1 u5_mult_82_S2_6_38 ( .A(u5_mult_82_ab_6__38_), .B(
        u5_mult_82_CARRYB_5__38_), .CI(u5_mult_82_SUMB_5__39_), .CO(
        u5_mult_82_CARRYB_6__38_), .S(u5_mult_82_SUMB_6__38_) );
  FA_X1 u5_mult_82_S2_6_37 ( .A(u5_mult_82_ab_6__37_), .B(
        u5_mult_82_CARRYB_5__37_), .CI(u5_mult_82_SUMB_5__38_), .CO(
        u5_mult_82_CARRYB_6__37_), .S(u5_mult_82_SUMB_6__37_) );
  FA_X1 u5_mult_82_S2_6_36 ( .A(u5_mult_82_ab_6__36_), .B(
        u5_mult_82_CARRYB_5__36_), .CI(u5_mult_82_SUMB_5__37_), .CO(
        u5_mult_82_CARRYB_6__36_), .S(u5_mult_82_SUMB_6__36_) );
  FA_X1 u5_mult_82_S2_6_35 ( .A(u5_mult_82_ab_6__35_), .B(
        u5_mult_82_CARRYB_5__35_), .CI(u5_mult_82_SUMB_5__36_), .CO(
        u5_mult_82_CARRYB_6__35_), .S(u5_mult_82_SUMB_6__35_) );
  FA_X1 u5_mult_82_S2_6_34 ( .A(u5_mult_82_ab_6__34_), .B(
        u5_mult_82_CARRYB_5__34_), .CI(u5_mult_82_SUMB_5__35_), .CO(
        u5_mult_82_CARRYB_6__34_), .S(u5_mult_82_SUMB_6__34_) );
  FA_X1 u5_mult_82_S2_6_33 ( .A(u5_mult_82_ab_6__33_), .B(
        u5_mult_82_CARRYB_5__33_), .CI(u5_mult_82_SUMB_5__34_), .CO(
        u5_mult_82_CARRYB_6__33_), .S(u5_mult_82_SUMB_6__33_) );
  FA_X1 u5_mult_82_S2_6_32 ( .A(u5_mult_82_ab_6__32_), .B(
        u5_mult_82_CARRYB_5__32_), .CI(u5_mult_82_SUMB_5__33_), .CO(
        u5_mult_82_CARRYB_6__32_), .S(u5_mult_82_SUMB_6__32_) );
  FA_X1 u5_mult_82_S2_6_31 ( .A(u5_mult_82_ab_6__31_), .B(
        u5_mult_82_CARRYB_5__31_), .CI(u5_mult_82_SUMB_5__32_), .CO(
        u5_mult_82_CARRYB_6__31_), .S(u5_mult_82_SUMB_6__31_) );
  FA_X1 u5_mult_82_S2_6_30 ( .A(u5_mult_82_ab_6__30_), .B(
        u5_mult_82_CARRYB_5__30_), .CI(u5_mult_82_SUMB_5__31_), .CO(
        u5_mult_82_CARRYB_6__30_), .S(u5_mult_82_SUMB_6__30_) );
  FA_X1 u5_mult_82_S2_6_29 ( .A(u5_mult_82_ab_6__29_), .B(
        u5_mult_82_CARRYB_5__29_), .CI(u5_mult_82_SUMB_5__30_), .CO(
        u5_mult_82_CARRYB_6__29_), .S(u5_mult_82_SUMB_6__29_) );
  FA_X1 u5_mult_82_S2_6_28 ( .A(u5_mult_82_ab_6__28_), .B(
        u5_mult_82_CARRYB_5__28_), .CI(u5_mult_82_SUMB_5__29_), .CO(
        u5_mult_82_CARRYB_6__28_), .S(u5_mult_82_SUMB_6__28_) );
  FA_X1 u5_mult_82_S2_6_27 ( .A(u5_mult_82_ab_6__27_), .B(
        u5_mult_82_CARRYB_5__27_), .CI(u5_mult_82_SUMB_5__28_), .CO(
        u5_mult_82_CARRYB_6__27_), .S(u5_mult_82_SUMB_6__27_) );
  FA_X1 u5_mult_82_S2_6_26 ( .A(u5_mult_82_ab_6__26_), .B(
        u5_mult_82_CARRYB_5__26_), .CI(u5_mult_82_SUMB_5__27_), .CO(
        u5_mult_82_CARRYB_6__26_), .S(u5_mult_82_SUMB_6__26_) );
  FA_X1 u5_mult_82_S2_6_25 ( .A(u5_mult_82_ab_6__25_), .B(
        u5_mult_82_CARRYB_5__25_), .CI(u5_mult_82_SUMB_5__26_), .CO(
        u5_mult_82_CARRYB_6__25_), .S(u5_mult_82_SUMB_6__25_) );
  FA_X1 u5_mult_82_S2_6_24 ( .A(u5_mult_82_ab_6__24_), .B(
        u5_mult_82_CARRYB_5__24_), .CI(u5_mult_82_SUMB_5__25_), .CO(
        u5_mult_82_CARRYB_6__24_), .S(u5_mult_82_SUMB_6__24_) );
  FA_X1 u5_mult_82_S2_6_23 ( .A(u5_mult_82_ab_6__23_), .B(
        u5_mult_82_CARRYB_5__23_), .CI(u5_mult_82_SUMB_5__24_), .CO(
        u5_mult_82_CARRYB_6__23_), .S(u5_mult_82_SUMB_6__23_) );
  FA_X1 u5_mult_82_S2_6_22 ( .A(u5_mult_82_ab_6__22_), .B(
        u5_mult_82_CARRYB_5__22_), .CI(u5_mult_82_SUMB_5__23_), .CO(
        u5_mult_82_CARRYB_6__22_), .S(u5_mult_82_SUMB_6__22_) );
  FA_X1 u5_mult_82_S2_6_21 ( .A(u5_mult_82_ab_6__21_), .B(
        u5_mult_82_CARRYB_5__21_), .CI(u5_mult_82_SUMB_5__22_), .CO(
        u5_mult_82_CARRYB_6__21_), .S(u5_mult_82_SUMB_6__21_) );
  FA_X1 u5_mult_82_S2_6_20 ( .A(u5_mult_82_ab_6__20_), .B(
        u5_mult_82_CARRYB_5__20_), .CI(u5_mult_82_SUMB_5__21_), .CO(
        u5_mult_82_CARRYB_6__20_), .S(u5_mult_82_SUMB_6__20_) );
  FA_X1 u5_mult_82_S2_6_19 ( .A(u5_mult_82_ab_6__19_), .B(
        u5_mult_82_CARRYB_5__19_), .CI(u5_mult_82_SUMB_5__20_), .CO(
        u5_mult_82_CARRYB_6__19_), .S(u5_mult_82_SUMB_6__19_) );
  FA_X1 u5_mult_82_S2_6_18 ( .A(u5_mult_82_ab_6__18_), .B(
        u5_mult_82_CARRYB_5__18_), .CI(u5_mult_82_SUMB_5__19_), .CO(
        u5_mult_82_CARRYB_6__18_), .S(u5_mult_82_SUMB_6__18_) );
  FA_X1 u5_mult_82_S2_6_17 ( .A(u5_mult_82_ab_6__17_), .B(
        u5_mult_82_CARRYB_5__17_), .CI(u5_mult_82_SUMB_5__18_), .CO(
        u5_mult_82_CARRYB_6__17_), .S(u5_mult_82_SUMB_6__17_) );
  FA_X1 u5_mult_82_S2_6_16 ( .A(u5_mult_82_ab_6__16_), .B(
        u5_mult_82_CARRYB_5__16_), .CI(u5_mult_82_SUMB_5__17_), .CO(
        u5_mult_82_CARRYB_6__16_), .S(u5_mult_82_SUMB_6__16_) );
  FA_X1 u5_mult_82_S2_6_15 ( .A(u5_mult_82_ab_6__15_), .B(
        u5_mult_82_CARRYB_5__15_), .CI(u5_mult_82_SUMB_5__16_), .CO(
        u5_mult_82_CARRYB_6__15_), .S(u5_mult_82_SUMB_6__15_) );
  FA_X1 u5_mult_82_S2_6_14 ( .A(u5_mult_82_ab_6__14_), .B(
        u5_mult_82_CARRYB_5__14_), .CI(u5_mult_82_SUMB_5__15_), .CO(
        u5_mult_82_CARRYB_6__14_), .S(u5_mult_82_SUMB_6__14_) );
  FA_X1 u5_mult_82_S2_6_13 ( .A(u5_mult_82_ab_6__13_), .B(
        u5_mult_82_CARRYB_5__13_), .CI(u5_mult_82_SUMB_5__14_), .CO(
        u5_mult_82_CARRYB_6__13_), .S(u5_mult_82_SUMB_6__13_) );
  FA_X1 u5_mult_82_S2_6_12 ( .A(u5_mult_82_ab_6__12_), .B(
        u5_mult_82_CARRYB_5__12_), .CI(u5_mult_82_SUMB_5__13_), .CO(
        u5_mult_82_CARRYB_6__12_), .S(u5_mult_82_SUMB_6__12_) );
  FA_X1 u5_mult_82_S2_6_11 ( .A(u5_mult_82_ab_6__11_), .B(
        u5_mult_82_CARRYB_5__11_), .CI(u5_mult_82_SUMB_5__12_), .CO(
        u5_mult_82_CARRYB_6__11_), .S(u5_mult_82_SUMB_6__11_) );
  FA_X1 u5_mult_82_S2_6_10 ( .A(u5_mult_82_ab_6__10_), .B(
        u5_mult_82_CARRYB_5__10_), .CI(u5_mult_82_SUMB_5__11_), .CO(
        u5_mult_82_CARRYB_6__10_), .S(u5_mult_82_SUMB_6__10_) );
  FA_X1 u5_mult_82_S2_6_9 ( .A(u5_mult_82_ab_6__9_), .B(
        u5_mult_82_CARRYB_5__9_), .CI(u5_mult_82_SUMB_5__10_), .CO(
        u5_mult_82_CARRYB_6__9_), .S(u5_mult_82_SUMB_6__9_) );
  FA_X1 u5_mult_82_S2_6_8 ( .A(u5_mult_82_ab_6__8_), .B(
        u5_mult_82_CARRYB_5__8_), .CI(u5_mult_82_SUMB_5__9_), .CO(
        u5_mult_82_CARRYB_6__8_), .S(u5_mult_82_SUMB_6__8_) );
  FA_X1 u5_mult_82_S2_6_7 ( .A(u5_mult_82_ab_6__7_), .B(
        u5_mult_82_CARRYB_5__7_), .CI(u5_mult_82_SUMB_5__8_), .CO(
        u5_mult_82_CARRYB_6__7_), .S(u5_mult_82_SUMB_6__7_) );
  FA_X1 u5_mult_82_S2_6_6 ( .A(u5_mult_82_ab_6__6_), .B(
        u5_mult_82_CARRYB_5__6_), .CI(u5_mult_82_SUMB_5__7_), .CO(
        u5_mult_82_CARRYB_6__6_), .S(u5_mult_82_SUMB_6__6_) );
  FA_X1 u5_mult_82_S2_6_5 ( .A(u5_mult_82_ab_6__5_), .B(
        u5_mult_82_CARRYB_5__5_), .CI(u5_mult_82_SUMB_5__6_), .CO(
        u5_mult_82_CARRYB_6__5_), .S(u5_mult_82_SUMB_6__5_) );
  FA_X1 u5_mult_82_S2_6_4 ( .A(u5_mult_82_ab_6__4_), .B(
        u5_mult_82_CARRYB_5__4_), .CI(u5_mult_82_SUMB_5__5_), .CO(
        u5_mult_82_CARRYB_6__4_), .S(u5_mult_82_SUMB_6__4_) );
  FA_X1 u5_mult_82_S2_6_3 ( .A(u5_mult_82_ab_6__3_), .B(
        u5_mult_82_CARRYB_5__3_), .CI(u5_mult_82_SUMB_5__4_), .CO(
        u5_mult_82_CARRYB_6__3_), .S(u5_mult_82_SUMB_6__3_) );
  FA_X1 u5_mult_82_S2_6_2 ( .A(u5_mult_82_ab_6__2_), .B(
        u5_mult_82_CARRYB_5__2_), .CI(u5_mult_82_SUMB_5__3_), .CO(
        u5_mult_82_CARRYB_6__2_), .S(u5_mult_82_SUMB_6__2_) );
  FA_X1 u5_mult_82_S2_6_1 ( .A(u5_mult_82_ab_6__1_), .B(
        u5_mult_82_CARRYB_5__1_), .CI(u5_mult_82_SUMB_5__2_), .CO(
        u5_mult_82_CARRYB_6__1_), .S(u5_mult_82_SUMB_6__1_) );
  FA_X1 u5_mult_82_S1_6_0 ( .A(u5_mult_82_ab_6__0_), .B(
        u5_mult_82_CARRYB_5__0_), .CI(u5_mult_82_SUMB_5__1_), .CO(
        u5_mult_82_CARRYB_6__0_), .S(u5_N6) );
  FA_X1 u5_mult_82_S3_7_51 ( .A(u5_mult_82_ab_7__51_), .B(
        u5_mult_82_CARRYB_6__51_), .CI(u5_mult_82_ab_6__52_), .CO(
        u5_mult_82_CARRYB_7__51_), .S(u5_mult_82_SUMB_7__51_) );
  FA_X1 u5_mult_82_S2_7_50 ( .A(u5_mult_82_ab_7__50_), .B(
        u5_mult_82_CARRYB_6__50_), .CI(u5_mult_82_SUMB_6__51_), .CO(
        u5_mult_82_CARRYB_7__50_), .S(u5_mult_82_SUMB_7__50_) );
  FA_X1 u5_mult_82_S2_7_49 ( .A(u5_mult_82_ab_7__49_), .B(
        u5_mult_82_CARRYB_6__49_), .CI(u5_mult_82_SUMB_6__50_), .CO(
        u5_mult_82_CARRYB_7__49_), .S(u5_mult_82_SUMB_7__49_) );
  FA_X1 u5_mult_82_S2_7_48 ( .A(u5_mult_82_ab_7__48_), .B(
        u5_mult_82_CARRYB_6__48_), .CI(u5_mult_82_SUMB_6__49_), .CO(
        u5_mult_82_CARRYB_7__48_), .S(u5_mult_82_SUMB_7__48_) );
  FA_X1 u5_mult_82_S2_7_47 ( .A(u5_mult_82_ab_7__47_), .B(
        u5_mult_82_CARRYB_6__47_), .CI(u5_mult_82_SUMB_6__48_), .CO(
        u5_mult_82_CARRYB_7__47_), .S(u5_mult_82_SUMB_7__47_) );
  FA_X1 u5_mult_82_S2_7_46 ( .A(u5_mult_82_ab_7__46_), .B(
        u5_mult_82_CARRYB_6__46_), .CI(u5_mult_82_SUMB_6__47_), .CO(
        u5_mult_82_CARRYB_7__46_), .S(u5_mult_82_SUMB_7__46_) );
  FA_X1 u5_mult_82_S2_7_45 ( .A(u5_mult_82_ab_7__45_), .B(
        u5_mult_82_CARRYB_6__45_), .CI(u5_mult_82_SUMB_6__46_), .CO(
        u5_mult_82_CARRYB_7__45_), .S(u5_mult_82_SUMB_7__45_) );
  FA_X1 u5_mult_82_S2_7_44 ( .A(u5_mult_82_ab_7__44_), .B(
        u5_mult_82_CARRYB_6__44_), .CI(u5_mult_82_SUMB_6__45_), .CO(
        u5_mult_82_CARRYB_7__44_), .S(u5_mult_82_SUMB_7__44_) );
  FA_X1 u5_mult_82_S2_7_43 ( .A(u5_mult_82_ab_7__43_), .B(
        u5_mult_82_CARRYB_6__43_), .CI(u5_mult_82_SUMB_6__44_), .CO(
        u5_mult_82_CARRYB_7__43_), .S(u5_mult_82_SUMB_7__43_) );
  FA_X1 u5_mult_82_S2_7_42 ( .A(u5_mult_82_ab_7__42_), .B(
        u5_mult_82_CARRYB_6__42_), .CI(u5_mult_82_SUMB_6__43_), .CO(
        u5_mult_82_CARRYB_7__42_), .S(u5_mult_82_SUMB_7__42_) );
  FA_X1 u5_mult_82_S2_7_41 ( .A(u5_mult_82_ab_7__41_), .B(
        u5_mult_82_CARRYB_6__41_), .CI(u5_mult_82_SUMB_6__42_), .CO(
        u5_mult_82_CARRYB_7__41_), .S(u5_mult_82_SUMB_7__41_) );
  FA_X1 u5_mult_82_S2_7_40 ( .A(u5_mult_82_ab_7__40_), .B(
        u5_mult_82_CARRYB_6__40_), .CI(u5_mult_82_SUMB_6__41_), .CO(
        u5_mult_82_CARRYB_7__40_), .S(u5_mult_82_SUMB_7__40_) );
  FA_X1 u5_mult_82_S2_7_39 ( .A(u5_mult_82_ab_7__39_), .B(
        u5_mult_82_CARRYB_6__39_), .CI(u5_mult_82_SUMB_6__40_), .CO(
        u5_mult_82_CARRYB_7__39_), .S(u5_mult_82_SUMB_7__39_) );
  FA_X1 u5_mult_82_S2_7_38 ( .A(u5_mult_82_ab_7__38_), .B(
        u5_mult_82_CARRYB_6__38_), .CI(u5_mult_82_SUMB_6__39_), .CO(
        u5_mult_82_CARRYB_7__38_), .S(u5_mult_82_SUMB_7__38_) );
  FA_X1 u5_mult_82_S2_7_37 ( .A(u5_mult_82_ab_7__37_), .B(
        u5_mult_82_CARRYB_6__37_), .CI(u5_mult_82_SUMB_6__38_), .CO(
        u5_mult_82_CARRYB_7__37_), .S(u5_mult_82_SUMB_7__37_) );
  FA_X1 u5_mult_82_S2_7_36 ( .A(u5_mult_82_ab_7__36_), .B(
        u5_mult_82_CARRYB_6__36_), .CI(u5_mult_82_SUMB_6__37_), .CO(
        u5_mult_82_CARRYB_7__36_), .S(u5_mult_82_SUMB_7__36_) );
  FA_X1 u5_mult_82_S2_7_35 ( .A(u5_mult_82_ab_7__35_), .B(
        u5_mult_82_CARRYB_6__35_), .CI(u5_mult_82_SUMB_6__36_), .CO(
        u5_mult_82_CARRYB_7__35_), .S(u5_mult_82_SUMB_7__35_) );
  FA_X1 u5_mult_82_S2_7_34 ( .A(u5_mult_82_ab_7__34_), .B(
        u5_mult_82_CARRYB_6__34_), .CI(u5_mult_82_SUMB_6__35_), .CO(
        u5_mult_82_CARRYB_7__34_), .S(u5_mult_82_SUMB_7__34_) );
  FA_X1 u5_mult_82_S2_7_33 ( .A(u5_mult_82_ab_7__33_), .B(
        u5_mult_82_CARRYB_6__33_), .CI(u5_mult_82_SUMB_6__34_), .CO(
        u5_mult_82_CARRYB_7__33_), .S(u5_mult_82_SUMB_7__33_) );
  FA_X1 u5_mult_82_S2_7_32 ( .A(u5_mult_82_ab_7__32_), .B(
        u5_mult_82_CARRYB_6__32_), .CI(u5_mult_82_SUMB_6__33_), .CO(
        u5_mult_82_CARRYB_7__32_), .S(u5_mult_82_SUMB_7__32_) );
  FA_X1 u5_mult_82_S2_7_31 ( .A(u5_mult_82_ab_7__31_), .B(
        u5_mult_82_CARRYB_6__31_), .CI(u5_mult_82_SUMB_6__32_), .CO(
        u5_mult_82_CARRYB_7__31_), .S(u5_mult_82_SUMB_7__31_) );
  FA_X1 u5_mult_82_S2_7_30 ( .A(u5_mult_82_ab_7__30_), .B(
        u5_mult_82_CARRYB_6__30_), .CI(u5_mult_82_SUMB_6__31_), .CO(
        u5_mult_82_CARRYB_7__30_), .S(u5_mult_82_SUMB_7__30_) );
  FA_X1 u5_mult_82_S2_7_29 ( .A(u5_mult_82_ab_7__29_), .B(
        u5_mult_82_CARRYB_6__29_), .CI(u5_mult_82_SUMB_6__30_), .CO(
        u5_mult_82_CARRYB_7__29_), .S(u5_mult_82_SUMB_7__29_) );
  FA_X1 u5_mult_82_S2_7_28 ( .A(u5_mult_82_ab_7__28_), .B(
        u5_mult_82_CARRYB_6__28_), .CI(u5_mult_82_SUMB_6__29_), .CO(
        u5_mult_82_CARRYB_7__28_), .S(u5_mult_82_SUMB_7__28_) );
  FA_X1 u5_mult_82_S2_7_27 ( .A(u5_mult_82_ab_7__27_), .B(
        u5_mult_82_CARRYB_6__27_), .CI(u5_mult_82_SUMB_6__28_), .CO(
        u5_mult_82_CARRYB_7__27_), .S(u5_mult_82_SUMB_7__27_) );
  FA_X1 u5_mult_82_S2_7_26 ( .A(u5_mult_82_ab_7__26_), .B(
        u5_mult_82_CARRYB_6__26_), .CI(u5_mult_82_SUMB_6__27_), .CO(
        u5_mult_82_CARRYB_7__26_), .S(u5_mult_82_SUMB_7__26_) );
  FA_X1 u5_mult_82_S2_7_25 ( .A(u5_mult_82_ab_7__25_), .B(
        u5_mult_82_CARRYB_6__25_), .CI(u5_mult_82_SUMB_6__26_), .CO(
        u5_mult_82_CARRYB_7__25_), .S(u5_mult_82_SUMB_7__25_) );
  FA_X1 u5_mult_82_S2_7_24 ( .A(u5_mult_82_ab_7__24_), .B(
        u5_mult_82_CARRYB_6__24_), .CI(u5_mult_82_SUMB_6__25_), .CO(
        u5_mult_82_CARRYB_7__24_), .S(u5_mult_82_SUMB_7__24_) );
  FA_X1 u5_mult_82_S2_7_23 ( .A(u5_mult_82_ab_7__23_), .B(
        u5_mult_82_CARRYB_6__23_), .CI(u5_mult_82_SUMB_6__24_), .CO(
        u5_mult_82_CARRYB_7__23_), .S(u5_mult_82_SUMB_7__23_) );
  FA_X1 u5_mult_82_S2_7_22 ( .A(u5_mult_82_ab_7__22_), .B(
        u5_mult_82_CARRYB_6__22_), .CI(u5_mult_82_SUMB_6__23_), .CO(
        u5_mult_82_CARRYB_7__22_), .S(u5_mult_82_SUMB_7__22_) );
  FA_X1 u5_mult_82_S2_7_21 ( .A(u5_mult_82_ab_7__21_), .B(
        u5_mult_82_CARRYB_6__21_), .CI(u5_mult_82_SUMB_6__22_), .CO(
        u5_mult_82_CARRYB_7__21_), .S(u5_mult_82_SUMB_7__21_) );
  FA_X1 u5_mult_82_S2_7_20 ( .A(u5_mult_82_ab_7__20_), .B(
        u5_mult_82_CARRYB_6__20_), .CI(u5_mult_82_SUMB_6__21_), .CO(
        u5_mult_82_CARRYB_7__20_), .S(u5_mult_82_SUMB_7__20_) );
  FA_X1 u5_mult_82_S2_7_19 ( .A(u5_mult_82_ab_7__19_), .B(
        u5_mult_82_CARRYB_6__19_), .CI(u5_mult_82_SUMB_6__20_), .CO(
        u5_mult_82_CARRYB_7__19_), .S(u5_mult_82_SUMB_7__19_) );
  FA_X1 u5_mult_82_S2_7_18 ( .A(u5_mult_82_ab_7__18_), .B(
        u5_mult_82_CARRYB_6__18_), .CI(u5_mult_82_SUMB_6__19_), .CO(
        u5_mult_82_CARRYB_7__18_), .S(u5_mult_82_SUMB_7__18_) );
  FA_X1 u5_mult_82_S2_7_17 ( .A(u5_mult_82_ab_7__17_), .B(
        u5_mult_82_CARRYB_6__17_), .CI(u5_mult_82_SUMB_6__18_), .CO(
        u5_mult_82_CARRYB_7__17_), .S(u5_mult_82_SUMB_7__17_) );
  FA_X1 u5_mult_82_S2_7_16 ( .A(u5_mult_82_ab_7__16_), .B(
        u5_mult_82_CARRYB_6__16_), .CI(u5_mult_82_SUMB_6__17_), .CO(
        u5_mult_82_CARRYB_7__16_), .S(u5_mult_82_SUMB_7__16_) );
  FA_X1 u5_mult_82_S2_7_15 ( .A(u5_mult_82_ab_7__15_), .B(
        u5_mult_82_CARRYB_6__15_), .CI(u5_mult_82_SUMB_6__16_), .CO(
        u5_mult_82_CARRYB_7__15_), .S(u5_mult_82_SUMB_7__15_) );
  FA_X1 u5_mult_82_S2_7_14 ( .A(u5_mult_82_ab_7__14_), .B(
        u5_mult_82_CARRYB_6__14_), .CI(u5_mult_82_SUMB_6__15_), .CO(
        u5_mult_82_CARRYB_7__14_), .S(u5_mult_82_SUMB_7__14_) );
  FA_X1 u5_mult_82_S2_7_13 ( .A(u5_mult_82_ab_7__13_), .B(
        u5_mult_82_CARRYB_6__13_), .CI(u5_mult_82_SUMB_6__14_), .CO(
        u5_mult_82_CARRYB_7__13_), .S(u5_mult_82_SUMB_7__13_) );
  FA_X1 u5_mult_82_S2_7_12 ( .A(u5_mult_82_ab_7__12_), .B(
        u5_mult_82_CARRYB_6__12_), .CI(u5_mult_82_SUMB_6__13_), .CO(
        u5_mult_82_CARRYB_7__12_), .S(u5_mult_82_SUMB_7__12_) );
  FA_X1 u5_mult_82_S2_7_11 ( .A(u5_mult_82_ab_7__11_), .B(
        u5_mult_82_CARRYB_6__11_), .CI(u5_mult_82_SUMB_6__12_), .CO(
        u5_mult_82_CARRYB_7__11_), .S(u5_mult_82_SUMB_7__11_) );
  FA_X1 u5_mult_82_S2_7_10 ( .A(u5_mult_82_ab_7__10_), .B(
        u5_mult_82_CARRYB_6__10_), .CI(u5_mult_82_SUMB_6__11_), .CO(
        u5_mult_82_CARRYB_7__10_), .S(u5_mult_82_SUMB_7__10_) );
  FA_X1 u5_mult_82_S2_7_9 ( .A(u5_mult_82_ab_7__9_), .B(
        u5_mult_82_CARRYB_6__9_), .CI(u5_mult_82_SUMB_6__10_), .CO(
        u5_mult_82_CARRYB_7__9_), .S(u5_mult_82_SUMB_7__9_) );
  FA_X1 u5_mult_82_S2_7_8 ( .A(u5_mult_82_ab_7__8_), .B(
        u5_mult_82_CARRYB_6__8_), .CI(u5_mult_82_SUMB_6__9_), .CO(
        u5_mult_82_CARRYB_7__8_), .S(u5_mult_82_SUMB_7__8_) );
  FA_X1 u5_mult_82_S2_7_7 ( .A(u5_mult_82_ab_7__7_), .B(
        u5_mult_82_CARRYB_6__7_), .CI(u5_mult_82_SUMB_6__8_), .CO(
        u5_mult_82_CARRYB_7__7_), .S(u5_mult_82_SUMB_7__7_) );
  FA_X1 u5_mult_82_S2_7_6 ( .A(u5_mult_82_ab_7__6_), .B(
        u5_mult_82_CARRYB_6__6_), .CI(u5_mult_82_SUMB_6__7_), .CO(
        u5_mult_82_CARRYB_7__6_), .S(u5_mult_82_SUMB_7__6_) );
  FA_X1 u5_mult_82_S2_7_5 ( .A(u5_mult_82_ab_7__5_), .B(
        u5_mult_82_CARRYB_6__5_), .CI(u5_mult_82_SUMB_6__6_), .CO(
        u5_mult_82_CARRYB_7__5_), .S(u5_mult_82_SUMB_7__5_) );
  FA_X1 u5_mult_82_S2_7_4 ( .A(u5_mult_82_ab_7__4_), .B(
        u5_mult_82_CARRYB_6__4_), .CI(u5_mult_82_SUMB_6__5_), .CO(
        u5_mult_82_CARRYB_7__4_), .S(u5_mult_82_SUMB_7__4_) );
  FA_X1 u5_mult_82_S2_7_3 ( .A(u5_mult_82_ab_7__3_), .B(
        u5_mult_82_CARRYB_6__3_), .CI(u5_mult_82_SUMB_6__4_), .CO(
        u5_mult_82_CARRYB_7__3_), .S(u5_mult_82_SUMB_7__3_) );
  FA_X1 u5_mult_82_S2_7_2 ( .A(u5_mult_82_ab_7__2_), .B(
        u5_mult_82_CARRYB_6__2_), .CI(u5_mult_82_SUMB_6__3_), .CO(
        u5_mult_82_CARRYB_7__2_), .S(u5_mult_82_SUMB_7__2_) );
  FA_X1 u5_mult_82_S2_7_1 ( .A(u5_mult_82_ab_7__1_), .B(
        u5_mult_82_CARRYB_6__1_), .CI(u5_mult_82_SUMB_6__2_), .CO(
        u5_mult_82_CARRYB_7__1_), .S(u5_mult_82_SUMB_7__1_) );
  FA_X1 u5_mult_82_S1_7_0 ( .A(u5_mult_82_ab_7__0_), .B(
        u5_mult_82_CARRYB_6__0_), .CI(u5_mult_82_SUMB_6__1_), .CO(
        u5_mult_82_CARRYB_7__0_), .S(u5_N7) );
  FA_X1 u5_mult_82_S3_8_51 ( .A(u5_mult_82_ab_8__51_), .B(
        u5_mult_82_CARRYB_7__51_), .CI(u5_mult_82_ab_7__52_), .CO(
        u5_mult_82_CARRYB_8__51_), .S(u5_mult_82_SUMB_8__51_) );
  FA_X1 u5_mult_82_S2_8_50 ( .A(u5_mult_82_ab_8__50_), .B(
        u5_mult_82_CARRYB_7__50_), .CI(u5_mult_82_SUMB_7__51_), .CO(
        u5_mult_82_CARRYB_8__50_), .S(u5_mult_82_SUMB_8__50_) );
  FA_X1 u5_mult_82_S2_8_49 ( .A(u5_mult_82_ab_8__49_), .B(
        u5_mult_82_CARRYB_7__49_), .CI(u5_mult_82_SUMB_7__50_), .CO(
        u5_mult_82_CARRYB_8__49_), .S(u5_mult_82_SUMB_8__49_) );
  FA_X1 u5_mult_82_S2_8_48 ( .A(u5_mult_82_ab_8__48_), .B(
        u5_mult_82_CARRYB_7__48_), .CI(u5_mult_82_SUMB_7__49_), .CO(
        u5_mult_82_CARRYB_8__48_), .S(u5_mult_82_SUMB_8__48_) );
  FA_X1 u5_mult_82_S2_8_47 ( .A(u5_mult_82_ab_8__47_), .B(
        u5_mult_82_CARRYB_7__47_), .CI(u5_mult_82_SUMB_7__48_), .CO(
        u5_mult_82_CARRYB_8__47_), .S(u5_mult_82_SUMB_8__47_) );
  FA_X1 u5_mult_82_S2_8_46 ( .A(u5_mult_82_ab_8__46_), .B(
        u5_mult_82_CARRYB_7__46_), .CI(u5_mult_82_SUMB_7__47_), .CO(
        u5_mult_82_CARRYB_8__46_), .S(u5_mult_82_SUMB_8__46_) );
  FA_X1 u5_mult_82_S2_8_45 ( .A(u5_mult_82_ab_8__45_), .B(
        u5_mult_82_CARRYB_7__45_), .CI(u5_mult_82_SUMB_7__46_), .CO(
        u5_mult_82_CARRYB_8__45_), .S(u5_mult_82_SUMB_8__45_) );
  FA_X1 u5_mult_82_S2_8_44 ( .A(u5_mult_82_ab_8__44_), .B(
        u5_mult_82_CARRYB_7__44_), .CI(u5_mult_82_SUMB_7__45_), .CO(
        u5_mult_82_CARRYB_8__44_), .S(u5_mult_82_SUMB_8__44_) );
  FA_X1 u5_mult_82_S2_8_43 ( .A(u5_mult_82_ab_8__43_), .B(
        u5_mult_82_CARRYB_7__43_), .CI(u5_mult_82_SUMB_7__44_), .CO(
        u5_mult_82_CARRYB_8__43_), .S(u5_mult_82_SUMB_8__43_) );
  FA_X1 u5_mult_82_S2_8_42 ( .A(u5_mult_82_ab_8__42_), .B(
        u5_mult_82_CARRYB_7__42_), .CI(u5_mult_82_SUMB_7__43_), .CO(
        u5_mult_82_CARRYB_8__42_), .S(u5_mult_82_SUMB_8__42_) );
  FA_X1 u5_mult_82_S2_8_41 ( .A(u5_mult_82_ab_8__41_), .B(
        u5_mult_82_CARRYB_7__41_), .CI(u5_mult_82_SUMB_7__42_), .CO(
        u5_mult_82_CARRYB_8__41_), .S(u5_mult_82_SUMB_8__41_) );
  FA_X1 u5_mult_82_S2_8_40 ( .A(u5_mult_82_ab_8__40_), .B(
        u5_mult_82_CARRYB_7__40_), .CI(u5_mult_82_SUMB_7__41_), .CO(
        u5_mult_82_CARRYB_8__40_), .S(u5_mult_82_SUMB_8__40_) );
  FA_X1 u5_mult_82_S2_8_39 ( .A(u5_mult_82_ab_8__39_), .B(
        u5_mult_82_CARRYB_7__39_), .CI(u5_mult_82_SUMB_7__40_), .CO(
        u5_mult_82_CARRYB_8__39_), .S(u5_mult_82_SUMB_8__39_) );
  FA_X1 u5_mult_82_S2_8_38 ( .A(u5_mult_82_ab_8__38_), .B(
        u5_mult_82_CARRYB_7__38_), .CI(u5_mult_82_SUMB_7__39_), .CO(
        u5_mult_82_CARRYB_8__38_), .S(u5_mult_82_SUMB_8__38_) );
  FA_X1 u5_mult_82_S2_8_37 ( .A(u5_mult_82_ab_8__37_), .B(
        u5_mult_82_CARRYB_7__37_), .CI(u5_mult_82_SUMB_7__38_), .CO(
        u5_mult_82_CARRYB_8__37_), .S(u5_mult_82_SUMB_8__37_) );
  FA_X1 u5_mult_82_S2_8_36 ( .A(u5_mult_82_ab_8__36_), .B(
        u5_mult_82_CARRYB_7__36_), .CI(u5_mult_82_SUMB_7__37_), .CO(
        u5_mult_82_CARRYB_8__36_), .S(u5_mult_82_SUMB_8__36_) );
  FA_X1 u5_mult_82_S2_8_35 ( .A(u5_mult_82_ab_8__35_), .B(
        u5_mult_82_CARRYB_7__35_), .CI(u5_mult_82_SUMB_7__36_), .CO(
        u5_mult_82_CARRYB_8__35_), .S(u5_mult_82_SUMB_8__35_) );
  FA_X1 u5_mult_82_S2_8_34 ( .A(u5_mult_82_ab_8__34_), .B(
        u5_mult_82_CARRYB_7__34_), .CI(u5_mult_82_SUMB_7__35_), .CO(
        u5_mult_82_CARRYB_8__34_), .S(u5_mult_82_SUMB_8__34_) );
  FA_X1 u5_mult_82_S2_8_33 ( .A(u5_mult_82_ab_8__33_), .B(
        u5_mult_82_CARRYB_7__33_), .CI(u5_mult_82_SUMB_7__34_), .CO(
        u5_mult_82_CARRYB_8__33_), .S(u5_mult_82_SUMB_8__33_) );
  FA_X1 u5_mult_82_S2_8_32 ( .A(u5_mult_82_ab_8__32_), .B(
        u5_mult_82_CARRYB_7__32_), .CI(u5_mult_82_SUMB_7__33_), .CO(
        u5_mult_82_CARRYB_8__32_), .S(u5_mult_82_SUMB_8__32_) );
  FA_X1 u5_mult_82_S2_8_31 ( .A(u5_mult_82_ab_8__31_), .B(
        u5_mult_82_CARRYB_7__31_), .CI(u5_mult_82_SUMB_7__32_), .CO(
        u5_mult_82_CARRYB_8__31_), .S(u5_mult_82_SUMB_8__31_) );
  FA_X1 u5_mult_82_S2_8_30 ( .A(u5_mult_82_ab_8__30_), .B(
        u5_mult_82_CARRYB_7__30_), .CI(u5_mult_82_SUMB_7__31_), .CO(
        u5_mult_82_CARRYB_8__30_), .S(u5_mult_82_SUMB_8__30_) );
  FA_X1 u5_mult_82_S2_8_29 ( .A(u5_mult_82_ab_8__29_), .B(
        u5_mult_82_CARRYB_7__29_), .CI(u5_mult_82_SUMB_7__30_), .CO(
        u5_mult_82_CARRYB_8__29_), .S(u5_mult_82_SUMB_8__29_) );
  FA_X1 u5_mult_82_S2_8_28 ( .A(u5_mult_82_ab_8__28_), .B(
        u5_mult_82_CARRYB_7__28_), .CI(u5_mult_82_SUMB_7__29_), .CO(
        u5_mult_82_CARRYB_8__28_), .S(u5_mult_82_SUMB_8__28_) );
  FA_X1 u5_mult_82_S2_8_27 ( .A(u5_mult_82_ab_8__27_), .B(
        u5_mult_82_CARRYB_7__27_), .CI(u5_mult_82_SUMB_7__28_), .CO(
        u5_mult_82_CARRYB_8__27_), .S(u5_mult_82_SUMB_8__27_) );
  FA_X1 u5_mult_82_S2_8_26 ( .A(u5_mult_82_ab_8__26_), .B(
        u5_mult_82_CARRYB_7__26_), .CI(u5_mult_82_SUMB_7__27_), .CO(
        u5_mult_82_CARRYB_8__26_), .S(u5_mult_82_SUMB_8__26_) );
  FA_X1 u5_mult_82_S2_8_25 ( .A(u5_mult_82_ab_8__25_), .B(
        u5_mult_82_CARRYB_7__25_), .CI(u5_mult_82_SUMB_7__26_), .CO(
        u5_mult_82_CARRYB_8__25_), .S(u5_mult_82_SUMB_8__25_) );
  FA_X1 u5_mult_82_S2_8_24 ( .A(u5_mult_82_ab_8__24_), .B(
        u5_mult_82_CARRYB_7__24_), .CI(u5_mult_82_SUMB_7__25_), .CO(
        u5_mult_82_CARRYB_8__24_), .S(u5_mult_82_SUMB_8__24_) );
  FA_X1 u5_mult_82_S2_8_23 ( .A(u5_mult_82_ab_8__23_), .B(
        u5_mult_82_CARRYB_7__23_), .CI(u5_mult_82_SUMB_7__24_), .CO(
        u5_mult_82_CARRYB_8__23_), .S(u5_mult_82_SUMB_8__23_) );
  FA_X1 u5_mult_82_S2_8_22 ( .A(u5_mult_82_ab_8__22_), .B(
        u5_mult_82_CARRYB_7__22_), .CI(u5_mult_82_SUMB_7__23_), .CO(
        u5_mult_82_CARRYB_8__22_), .S(u5_mult_82_SUMB_8__22_) );
  FA_X1 u5_mult_82_S2_8_21 ( .A(u5_mult_82_ab_8__21_), .B(
        u5_mult_82_CARRYB_7__21_), .CI(u5_mult_82_SUMB_7__22_), .CO(
        u5_mult_82_CARRYB_8__21_), .S(u5_mult_82_SUMB_8__21_) );
  FA_X1 u5_mult_82_S2_8_20 ( .A(u5_mult_82_ab_8__20_), .B(
        u5_mult_82_CARRYB_7__20_), .CI(u5_mult_82_SUMB_7__21_), .CO(
        u5_mult_82_CARRYB_8__20_), .S(u5_mult_82_SUMB_8__20_) );
  FA_X1 u5_mult_82_S2_8_19 ( .A(u5_mult_82_ab_8__19_), .B(
        u5_mult_82_CARRYB_7__19_), .CI(u5_mult_82_SUMB_7__20_), .CO(
        u5_mult_82_CARRYB_8__19_), .S(u5_mult_82_SUMB_8__19_) );
  FA_X1 u5_mult_82_S2_8_18 ( .A(u5_mult_82_ab_8__18_), .B(
        u5_mult_82_CARRYB_7__18_), .CI(u5_mult_82_SUMB_7__19_), .CO(
        u5_mult_82_CARRYB_8__18_), .S(u5_mult_82_SUMB_8__18_) );
  FA_X1 u5_mult_82_S2_8_17 ( .A(u5_mult_82_ab_8__17_), .B(
        u5_mult_82_CARRYB_7__17_), .CI(u5_mult_82_SUMB_7__18_), .CO(
        u5_mult_82_CARRYB_8__17_), .S(u5_mult_82_SUMB_8__17_) );
  FA_X1 u5_mult_82_S2_8_16 ( .A(u5_mult_82_ab_8__16_), .B(
        u5_mult_82_CARRYB_7__16_), .CI(u5_mult_82_SUMB_7__17_), .CO(
        u5_mult_82_CARRYB_8__16_), .S(u5_mult_82_SUMB_8__16_) );
  FA_X1 u5_mult_82_S2_8_15 ( .A(u5_mult_82_ab_8__15_), .B(
        u5_mult_82_CARRYB_7__15_), .CI(u5_mult_82_SUMB_7__16_), .CO(
        u5_mult_82_CARRYB_8__15_), .S(u5_mult_82_SUMB_8__15_) );
  FA_X1 u5_mult_82_S2_8_14 ( .A(u5_mult_82_ab_8__14_), .B(
        u5_mult_82_CARRYB_7__14_), .CI(u5_mult_82_SUMB_7__15_), .CO(
        u5_mult_82_CARRYB_8__14_), .S(u5_mult_82_SUMB_8__14_) );
  FA_X1 u5_mult_82_S2_8_13 ( .A(u5_mult_82_ab_8__13_), .B(
        u5_mult_82_CARRYB_7__13_), .CI(u5_mult_82_SUMB_7__14_), .CO(
        u5_mult_82_CARRYB_8__13_), .S(u5_mult_82_SUMB_8__13_) );
  FA_X1 u5_mult_82_S2_8_12 ( .A(u5_mult_82_ab_8__12_), .B(
        u5_mult_82_CARRYB_7__12_), .CI(u5_mult_82_SUMB_7__13_), .CO(
        u5_mult_82_CARRYB_8__12_), .S(u5_mult_82_SUMB_8__12_) );
  FA_X1 u5_mult_82_S2_8_11 ( .A(u5_mult_82_ab_8__11_), .B(
        u5_mult_82_CARRYB_7__11_), .CI(u5_mult_82_SUMB_7__12_), .CO(
        u5_mult_82_CARRYB_8__11_), .S(u5_mult_82_SUMB_8__11_) );
  FA_X1 u5_mult_82_S2_8_10 ( .A(u5_mult_82_ab_8__10_), .B(
        u5_mult_82_CARRYB_7__10_), .CI(u5_mult_82_SUMB_7__11_), .CO(
        u5_mult_82_CARRYB_8__10_), .S(u5_mult_82_SUMB_8__10_) );
  FA_X1 u5_mult_82_S2_8_9 ( .A(u5_mult_82_ab_8__9_), .B(
        u5_mult_82_CARRYB_7__9_), .CI(u5_mult_82_SUMB_7__10_), .CO(
        u5_mult_82_CARRYB_8__9_), .S(u5_mult_82_SUMB_8__9_) );
  FA_X1 u5_mult_82_S2_8_8 ( .A(u5_mult_82_ab_8__8_), .B(
        u5_mult_82_CARRYB_7__8_), .CI(u5_mult_82_SUMB_7__9_), .CO(
        u5_mult_82_CARRYB_8__8_), .S(u5_mult_82_SUMB_8__8_) );
  FA_X1 u5_mult_82_S2_8_7 ( .A(u5_mult_82_ab_8__7_), .B(
        u5_mult_82_CARRYB_7__7_), .CI(u5_mult_82_SUMB_7__8_), .CO(
        u5_mult_82_CARRYB_8__7_), .S(u5_mult_82_SUMB_8__7_) );
  FA_X1 u5_mult_82_S2_8_6 ( .A(u5_mult_82_ab_8__6_), .B(
        u5_mult_82_CARRYB_7__6_), .CI(u5_mult_82_SUMB_7__7_), .CO(
        u5_mult_82_CARRYB_8__6_), .S(u5_mult_82_SUMB_8__6_) );
  FA_X1 u5_mult_82_S2_8_5 ( .A(u5_mult_82_ab_8__5_), .B(
        u5_mult_82_CARRYB_7__5_), .CI(u5_mult_82_SUMB_7__6_), .CO(
        u5_mult_82_CARRYB_8__5_), .S(u5_mult_82_SUMB_8__5_) );
  FA_X1 u5_mult_82_S2_8_4 ( .A(u5_mult_82_ab_8__4_), .B(
        u5_mult_82_CARRYB_7__4_), .CI(u5_mult_82_SUMB_7__5_), .CO(
        u5_mult_82_CARRYB_8__4_), .S(u5_mult_82_SUMB_8__4_) );
  FA_X1 u5_mult_82_S2_8_3 ( .A(u5_mult_82_ab_8__3_), .B(
        u5_mult_82_CARRYB_7__3_), .CI(u5_mult_82_SUMB_7__4_), .CO(
        u5_mult_82_CARRYB_8__3_), .S(u5_mult_82_SUMB_8__3_) );
  FA_X1 u5_mult_82_S2_8_2 ( .A(u5_mult_82_ab_8__2_), .B(
        u5_mult_82_CARRYB_7__2_), .CI(u5_mult_82_SUMB_7__3_), .CO(
        u5_mult_82_CARRYB_8__2_), .S(u5_mult_82_SUMB_8__2_) );
  FA_X1 u5_mult_82_S2_8_1 ( .A(u5_mult_82_ab_8__1_), .B(
        u5_mult_82_CARRYB_7__1_), .CI(u5_mult_82_SUMB_7__2_), .CO(
        u5_mult_82_CARRYB_8__1_), .S(u5_mult_82_SUMB_8__1_) );
  FA_X1 u5_mult_82_S1_8_0 ( .A(u5_mult_82_ab_8__0_), .B(
        u5_mult_82_CARRYB_7__0_), .CI(u5_mult_82_SUMB_7__1_), .CO(
        u5_mult_82_CARRYB_8__0_), .S(u5_N8) );
  FA_X1 u5_mult_82_S3_9_51 ( .A(u5_mult_82_ab_9__51_), .B(
        u5_mult_82_CARRYB_8__51_), .CI(u5_mult_82_ab_8__52_), .CO(
        u5_mult_82_CARRYB_9__51_), .S(u5_mult_82_SUMB_9__51_) );
  FA_X1 u5_mult_82_S2_9_50 ( .A(u5_mult_82_ab_9__50_), .B(
        u5_mult_82_CARRYB_8__50_), .CI(u5_mult_82_SUMB_8__51_), .CO(
        u5_mult_82_CARRYB_9__50_), .S(u5_mult_82_SUMB_9__50_) );
  FA_X1 u5_mult_82_S2_9_49 ( .A(u5_mult_82_ab_9__49_), .B(
        u5_mult_82_CARRYB_8__49_), .CI(u5_mult_82_SUMB_8__50_), .CO(
        u5_mult_82_CARRYB_9__49_), .S(u5_mult_82_SUMB_9__49_) );
  FA_X1 u5_mult_82_S2_9_48 ( .A(u5_mult_82_ab_9__48_), .B(
        u5_mult_82_CARRYB_8__48_), .CI(u5_mult_82_SUMB_8__49_), .CO(
        u5_mult_82_CARRYB_9__48_), .S(u5_mult_82_SUMB_9__48_) );
  FA_X1 u5_mult_82_S2_9_47 ( .A(u5_mult_82_ab_9__47_), .B(
        u5_mult_82_CARRYB_8__47_), .CI(u5_mult_82_SUMB_8__48_), .CO(
        u5_mult_82_CARRYB_9__47_), .S(u5_mult_82_SUMB_9__47_) );
  FA_X1 u5_mult_82_S2_9_46 ( .A(u5_mult_82_ab_9__46_), .B(
        u5_mult_82_CARRYB_8__46_), .CI(u5_mult_82_SUMB_8__47_), .CO(
        u5_mult_82_CARRYB_9__46_), .S(u5_mult_82_SUMB_9__46_) );
  FA_X1 u5_mult_82_S2_9_45 ( .A(u5_mult_82_ab_9__45_), .B(
        u5_mult_82_CARRYB_8__45_), .CI(u5_mult_82_SUMB_8__46_), .CO(
        u5_mult_82_CARRYB_9__45_), .S(u5_mult_82_SUMB_9__45_) );
  FA_X1 u5_mult_82_S2_9_44 ( .A(u5_mult_82_ab_9__44_), .B(
        u5_mult_82_CARRYB_8__44_), .CI(u5_mult_82_SUMB_8__45_), .CO(
        u5_mult_82_CARRYB_9__44_), .S(u5_mult_82_SUMB_9__44_) );
  FA_X1 u5_mult_82_S2_9_43 ( .A(u5_mult_82_ab_9__43_), .B(
        u5_mult_82_CARRYB_8__43_), .CI(u5_mult_82_SUMB_8__44_), .CO(
        u5_mult_82_CARRYB_9__43_), .S(u5_mult_82_SUMB_9__43_) );
  FA_X1 u5_mult_82_S2_9_42 ( .A(u5_mult_82_ab_9__42_), .B(
        u5_mult_82_CARRYB_8__42_), .CI(u5_mult_82_SUMB_8__43_), .CO(
        u5_mult_82_CARRYB_9__42_), .S(u5_mult_82_SUMB_9__42_) );
  FA_X1 u5_mult_82_S2_9_41 ( .A(u5_mult_82_ab_9__41_), .B(
        u5_mult_82_CARRYB_8__41_), .CI(u5_mult_82_SUMB_8__42_), .CO(
        u5_mult_82_CARRYB_9__41_), .S(u5_mult_82_SUMB_9__41_) );
  FA_X1 u5_mult_82_S2_9_40 ( .A(u5_mult_82_ab_9__40_), .B(
        u5_mult_82_CARRYB_8__40_), .CI(u5_mult_82_SUMB_8__41_), .CO(
        u5_mult_82_CARRYB_9__40_), .S(u5_mult_82_SUMB_9__40_) );
  FA_X1 u5_mult_82_S2_9_39 ( .A(u5_mult_82_ab_9__39_), .B(
        u5_mult_82_CARRYB_8__39_), .CI(u5_mult_82_SUMB_8__40_), .CO(
        u5_mult_82_CARRYB_9__39_), .S(u5_mult_82_SUMB_9__39_) );
  FA_X1 u5_mult_82_S2_9_38 ( .A(u5_mult_82_ab_9__38_), .B(
        u5_mult_82_CARRYB_8__38_), .CI(u5_mult_82_SUMB_8__39_), .CO(
        u5_mult_82_CARRYB_9__38_), .S(u5_mult_82_SUMB_9__38_) );
  FA_X1 u5_mult_82_S2_9_37 ( .A(u5_mult_82_ab_9__37_), .B(
        u5_mult_82_CARRYB_8__37_), .CI(u5_mult_82_SUMB_8__38_), .CO(
        u5_mult_82_CARRYB_9__37_), .S(u5_mult_82_SUMB_9__37_) );
  FA_X1 u5_mult_82_S2_9_36 ( .A(u5_mult_82_ab_9__36_), .B(
        u5_mult_82_CARRYB_8__36_), .CI(u5_mult_82_SUMB_8__37_), .CO(
        u5_mult_82_CARRYB_9__36_), .S(u5_mult_82_SUMB_9__36_) );
  FA_X1 u5_mult_82_S2_9_35 ( .A(u5_mult_82_ab_9__35_), .B(
        u5_mult_82_CARRYB_8__35_), .CI(u5_mult_82_SUMB_8__36_), .CO(
        u5_mult_82_CARRYB_9__35_), .S(u5_mult_82_SUMB_9__35_) );
  FA_X1 u5_mult_82_S2_9_34 ( .A(u5_mult_82_ab_9__34_), .B(
        u5_mult_82_CARRYB_8__34_), .CI(u5_mult_82_SUMB_8__35_), .CO(
        u5_mult_82_CARRYB_9__34_), .S(u5_mult_82_SUMB_9__34_) );
  FA_X1 u5_mult_82_S2_9_33 ( .A(u5_mult_82_ab_9__33_), .B(
        u5_mult_82_CARRYB_8__33_), .CI(u5_mult_82_SUMB_8__34_), .CO(
        u5_mult_82_CARRYB_9__33_), .S(u5_mult_82_SUMB_9__33_) );
  FA_X1 u5_mult_82_S2_9_32 ( .A(u5_mult_82_ab_9__32_), .B(
        u5_mult_82_CARRYB_8__32_), .CI(u5_mult_82_SUMB_8__33_), .CO(
        u5_mult_82_CARRYB_9__32_), .S(u5_mult_82_SUMB_9__32_) );
  FA_X1 u5_mult_82_S2_9_31 ( .A(u5_mult_82_ab_9__31_), .B(
        u5_mult_82_CARRYB_8__31_), .CI(u5_mult_82_SUMB_8__32_), .CO(
        u5_mult_82_CARRYB_9__31_), .S(u5_mult_82_SUMB_9__31_) );
  FA_X1 u5_mult_82_S2_9_30 ( .A(u5_mult_82_ab_9__30_), .B(
        u5_mult_82_CARRYB_8__30_), .CI(u5_mult_82_SUMB_8__31_), .CO(
        u5_mult_82_CARRYB_9__30_), .S(u5_mult_82_SUMB_9__30_) );
  FA_X1 u5_mult_82_S2_9_29 ( .A(u5_mult_82_ab_9__29_), .B(
        u5_mult_82_CARRYB_8__29_), .CI(u5_mult_82_SUMB_8__30_), .CO(
        u5_mult_82_CARRYB_9__29_), .S(u5_mult_82_SUMB_9__29_) );
  FA_X1 u5_mult_82_S2_9_28 ( .A(u5_mult_82_ab_9__28_), .B(
        u5_mult_82_CARRYB_8__28_), .CI(u5_mult_82_SUMB_8__29_), .CO(
        u5_mult_82_CARRYB_9__28_), .S(u5_mult_82_SUMB_9__28_) );
  FA_X1 u5_mult_82_S2_9_27 ( .A(u5_mult_82_ab_9__27_), .B(
        u5_mult_82_CARRYB_8__27_), .CI(u5_mult_82_SUMB_8__28_), .CO(
        u5_mult_82_CARRYB_9__27_), .S(u5_mult_82_SUMB_9__27_) );
  FA_X1 u5_mult_82_S2_9_26 ( .A(u5_mult_82_ab_9__26_), .B(
        u5_mult_82_CARRYB_8__26_), .CI(u5_mult_82_SUMB_8__27_), .CO(
        u5_mult_82_CARRYB_9__26_), .S(u5_mult_82_SUMB_9__26_) );
  FA_X1 u5_mult_82_S2_9_25 ( .A(u5_mult_82_ab_9__25_), .B(
        u5_mult_82_CARRYB_8__25_), .CI(u5_mult_82_SUMB_8__26_), .CO(
        u5_mult_82_CARRYB_9__25_), .S(u5_mult_82_SUMB_9__25_) );
  FA_X1 u5_mult_82_S2_9_24 ( .A(u5_mult_82_ab_9__24_), .B(
        u5_mult_82_CARRYB_8__24_), .CI(u5_mult_82_SUMB_8__25_), .CO(
        u5_mult_82_CARRYB_9__24_), .S(u5_mult_82_SUMB_9__24_) );
  FA_X1 u5_mult_82_S2_9_23 ( .A(u5_mult_82_ab_9__23_), .B(
        u5_mult_82_CARRYB_8__23_), .CI(u5_mult_82_SUMB_8__24_), .CO(
        u5_mult_82_CARRYB_9__23_), .S(u5_mult_82_SUMB_9__23_) );
  FA_X1 u5_mult_82_S2_9_22 ( .A(u5_mult_82_ab_9__22_), .B(
        u5_mult_82_CARRYB_8__22_), .CI(u5_mult_82_SUMB_8__23_), .CO(
        u5_mult_82_CARRYB_9__22_), .S(u5_mult_82_SUMB_9__22_) );
  FA_X1 u5_mult_82_S2_9_21 ( .A(u5_mult_82_ab_9__21_), .B(
        u5_mult_82_CARRYB_8__21_), .CI(u5_mult_82_SUMB_8__22_), .CO(
        u5_mult_82_CARRYB_9__21_), .S(u5_mult_82_SUMB_9__21_) );
  FA_X1 u5_mult_82_S2_9_20 ( .A(u5_mult_82_ab_9__20_), .B(
        u5_mult_82_CARRYB_8__20_), .CI(u5_mult_82_SUMB_8__21_), .CO(
        u5_mult_82_CARRYB_9__20_), .S(u5_mult_82_SUMB_9__20_) );
  FA_X1 u5_mult_82_S2_9_19 ( .A(u5_mult_82_ab_9__19_), .B(
        u5_mult_82_CARRYB_8__19_), .CI(u5_mult_82_SUMB_8__20_), .CO(
        u5_mult_82_CARRYB_9__19_), .S(u5_mult_82_SUMB_9__19_) );
  FA_X1 u5_mult_82_S2_9_18 ( .A(u5_mult_82_ab_9__18_), .B(
        u5_mult_82_CARRYB_8__18_), .CI(u5_mult_82_SUMB_8__19_), .CO(
        u5_mult_82_CARRYB_9__18_), .S(u5_mult_82_SUMB_9__18_) );
  FA_X1 u5_mult_82_S2_9_17 ( .A(u5_mult_82_ab_9__17_), .B(
        u5_mult_82_CARRYB_8__17_), .CI(u5_mult_82_SUMB_8__18_), .CO(
        u5_mult_82_CARRYB_9__17_), .S(u5_mult_82_SUMB_9__17_) );
  FA_X1 u5_mult_82_S2_9_16 ( .A(u5_mult_82_ab_9__16_), .B(
        u5_mult_82_CARRYB_8__16_), .CI(u5_mult_82_SUMB_8__17_), .CO(
        u5_mult_82_CARRYB_9__16_), .S(u5_mult_82_SUMB_9__16_) );
  FA_X1 u5_mult_82_S2_9_15 ( .A(u5_mult_82_ab_9__15_), .B(
        u5_mult_82_CARRYB_8__15_), .CI(u5_mult_82_SUMB_8__16_), .CO(
        u5_mult_82_CARRYB_9__15_), .S(u5_mult_82_SUMB_9__15_) );
  FA_X1 u5_mult_82_S2_9_14 ( .A(u5_mult_82_ab_9__14_), .B(
        u5_mult_82_CARRYB_8__14_), .CI(u5_mult_82_SUMB_8__15_), .CO(
        u5_mult_82_CARRYB_9__14_), .S(u5_mult_82_SUMB_9__14_) );
  FA_X1 u5_mult_82_S2_9_13 ( .A(u5_mult_82_ab_9__13_), .B(
        u5_mult_82_CARRYB_8__13_), .CI(u5_mult_82_SUMB_8__14_), .CO(
        u5_mult_82_CARRYB_9__13_), .S(u5_mult_82_SUMB_9__13_) );
  FA_X1 u5_mult_82_S2_9_12 ( .A(u5_mult_82_ab_9__12_), .B(
        u5_mult_82_CARRYB_8__12_), .CI(u5_mult_82_SUMB_8__13_), .CO(
        u5_mult_82_CARRYB_9__12_), .S(u5_mult_82_SUMB_9__12_) );
  FA_X1 u5_mult_82_S2_9_11 ( .A(u5_mult_82_ab_9__11_), .B(
        u5_mult_82_CARRYB_8__11_), .CI(u5_mult_82_SUMB_8__12_), .CO(
        u5_mult_82_CARRYB_9__11_), .S(u5_mult_82_SUMB_9__11_) );
  FA_X1 u5_mult_82_S2_9_10 ( .A(u5_mult_82_ab_9__10_), .B(
        u5_mult_82_CARRYB_8__10_), .CI(u5_mult_82_SUMB_8__11_), .CO(
        u5_mult_82_CARRYB_9__10_), .S(u5_mult_82_SUMB_9__10_) );
  FA_X1 u5_mult_82_S2_9_9 ( .A(u5_mult_82_ab_9__9_), .B(
        u5_mult_82_CARRYB_8__9_), .CI(u5_mult_82_SUMB_8__10_), .CO(
        u5_mult_82_CARRYB_9__9_), .S(u5_mult_82_SUMB_9__9_) );
  FA_X1 u5_mult_82_S2_9_8 ( .A(u5_mult_82_ab_9__8_), .B(
        u5_mult_82_CARRYB_8__8_), .CI(u5_mult_82_SUMB_8__9_), .CO(
        u5_mult_82_CARRYB_9__8_), .S(u5_mult_82_SUMB_9__8_) );
  FA_X1 u5_mult_82_S2_9_7 ( .A(u5_mult_82_ab_9__7_), .B(
        u5_mult_82_CARRYB_8__7_), .CI(u5_mult_82_SUMB_8__8_), .CO(
        u5_mult_82_CARRYB_9__7_), .S(u5_mult_82_SUMB_9__7_) );
  FA_X1 u5_mult_82_S2_9_6 ( .A(u5_mult_82_ab_9__6_), .B(
        u5_mult_82_CARRYB_8__6_), .CI(u5_mult_82_SUMB_8__7_), .CO(
        u5_mult_82_CARRYB_9__6_), .S(u5_mult_82_SUMB_9__6_) );
  FA_X1 u5_mult_82_S2_9_5 ( .A(u5_mult_82_ab_9__5_), .B(
        u5_mult_82_CARRYB_8__5_), .CI(u5_mult_82_SUMB_8__6_), .CO(
        u5_mult_82_CARRYB_9__5_), .S(u5_mult_82_SUMB_9__5_) );
  FA_X1 u5_mult_82_S2_9_4 ( .A(u5_mult_82_ab_9__4_), .B(
        u5_mult_82_CARRYB_8__4_), .CI(u5_mult_82_SUMB_8__5_), .CO(
        u5_mult_82_CARRYB_9__4_), .S(u5_mult_82_SUMB_9__4_) );
  FA_X1 u5_mult_82_S2_9_3 ( .A(u5_mult_82_ab_9__3_), .B(
        u5_mult_82_CARRYB_8__3_), .CI(u5_mult_82_SUMB_8__4_), .CO(
        u5_mult_82_CARRYB_9__3_), .S(u5_mult_82_SUMB_9__3_) );
  FA_X1 u5_mult_82_S2_9_2 ( .A(u5_mult_82_ab_9__2_), .B(
        u5_mult_82_CARRYB_8__2_), .CI(u5_mult_82_SUMB_8__3_), .CO(
        u5_mult_82_CARRYB_9__2_), .S(u5_mult_82_SUMB_9__2_) );
  FA_X1 u5_mult_82_S2_9_1 ( .A(u5_mult_82_ab_9__1_), .B(
        u5_mult_82_CARRYB_8__1_), .CI(u5_mult_82_SUMB_8__2_), .CO(
        u5_mult_82_CARRYB_9__1_), .S(u5_mult_82_SUMB_9__1_) );
  FA_X1 u5_mult_82_S1_9_0 ( .A(u5_mult_82_ab_9__0_), .B(
        u5_mult_82_CARRYB_8__0_), .CI(u5_mult_82_SUMB_8__1_), .CO(
        u5_mult_82_CARRYB_9__0_), .S(u5_N9) );
  FA_X1 u5_mult_82_S3_10_51 ( .A(u5_mult_82_ab_10__51_), .B(
        u5_mult_82_CARRYB_9__51_), .CI(u5_mult_82_ab_9__52_), .CO(
        u5_mult_82_CARRYB_10__51_), .S(u5_mult_82_SUMB_10__51_) );
  FA_X1 u5_mult_82_S2_10_50 ( .A(u5_mult_82_ab_10__50_), .B(
        u5_mult_82_CARRYB_9__50_), .CI(u5_mult_82_SUMB_9__51_), .CO(
        u5_mult_82_CARRYB_10__50_), .S(u5_mult_82_SUMB_10__50_) );
  FA_X1 u5_mult_82_S2_10_49 ( .A(u5_mult_82_ab_10__49_), .B(
        u5_mult_82_CARRYB_9__49_), .CI(u5_mult_82_SUMB_9__50_), .CO(
        u5_mult_82_CARRYB_10__49_), .S(u5_mult_82_SUMB_10__49_) );
  FA_X1 u5_mult_82_S2_10_48 ( .A(u5_mult_82_ab_10__48_), .B(
        u5_mult_82_CARRYB_9__48_), .CI(u5_mult_82_SUMB_9__49_), .CO(
        u5_mult_82_CARRYB_10__48_), .S(u5_mult_82_SUMB_10__48_) );
  FA_X1 u5_mult_82_S2_10_47 ( .A(u5_mult_82_ab_10__47_), .B(
        u5_mult_82_CARRYB_9__47_), .CI(u5_mult_82_SUMB_9__48_), .CO(
        u5_mult_82_CARRYB_10__47_), .S(u5_mult_82_SUMB_10__47_) );
  FA_X1 u5_mult_82_S2_10_46 ( .A(u5_mult_82_ab_10__46_), .B(
        u5_mult_82_CARRYB_9__46_), .CI(u5_mult_82_SUMB_9__47_), .CO(
        u5_mult_82_CARRYB_10__46_), .S(u5_mult_82_SUMB_10__46_) );
  FA_X1 u5_mult_82_S2_10_45 ( .A(u5_mult_82_ab_10__45_), .B(
        u5_mult_82_CARRYB_9__45_), .CI(u5_mult_82_SUMB_9__46_), .CO(
        u5_mult_82_CARRYB_10__45_), .S(u5_mult_82_SUMB_10__45_) );
  FA_X1 u5_mult_82_S2_10_44 ( .A(u5_mult_82_ab_10__44_), .B(
        u5_mult_82_CARRYB_9__44_), .CI(u5_mult_82_SUMB_9__45_), .CO(
        u5_mult_82_CARRYB_10__44_), .S(u5_mult_82_SUMB_10__44_) );
  FA_X1 u5_mult_82_S2_10_43 ( .A(u5_mult_82_ab_10__43_), .B(
        u5_mult_82_CARRYB_9__43_), .CI(u5_mult_82_SUMB_9__44_), .CO(
        u5_mult_82_CARRYB_10__43_), .S(u5_mult_82_SUMB_10__43_) );
  FA_X1 u5_mult_82_S2_10_42 ( .A(u5_mult_82_ab_10__42_), .B(
        u5_mult_82_CARRYB_9__42_), .CI(u5_mult_82_SUMB_9__43_), .CO(
        u5_mult_82_CARRYB_10__42_), .S(u5_mult_82_SUMB_10__42_) );
  FA_X1 u5_mult_82_S2_10_41 ( .A(u5_mult_82_ab_10__41_), .B(
        u5_mult_82_CARRYB_9__41_), .CI(u5_mult_82_SUMB_9__42_), .CO(
        u5_mult_82_CARRYB_10__41_), .S(u5_mult_82_SUMB_10__41_) );
  FA_X1 u5_mult_82_S2_10_40 ( .A(u5_mult_82_ab_10__40_), .B(
        u5_mult_82_CARRYB_9__40_), .CI(u5_mult_82_SUMB_9__41_), .CO(
        u5_mult_82_CARRYB_10__40_), .S(u5_mult_82_SUMB_10__40_) );
  FA_X1 u5_mult_82_S2_10_39 ( .A(u5_mult_82_ab_10__39_), .B(
        u5_mult_82_CARRYB_9__39_), .CI(u5_mult_82_SUMB_9__40_), .CO(
        u5_mult_82_CARRYB_10__39_), .S(u5_mult_82_SUMB_10__39_) );
  FA_X1 u5_mult_82_S2_10_38 ( .A(u5_mult_82_ab_10__38_), .B(
        u5_mult_82_CARRYB_9__38_), .CI(u5_mult_82_SUMB_9__39_), .CO(
        u5_mult_82_CARRYB_10__38_), .S(u5_mult_82_SUMB_10__38_) );
  FA_X1 u5_mult_82_S2_10_37 ( .A(u5_mult_82_ab_10__37_), .B(
        u5_mult_82_CARRYB_9__37_), .CI(u5_mult_82_SUMB_9__38_), .CO(
        u5_mult_82_CARRYB_10__37_), .S(u5_mult_82_SUMB_10__37_) );
  FA_X1 u5_mult_82_S2_10_36 ( .A(u5_mult_82_ab_10__36_), .B(
        u5_mult_82_CARRYB_9__36_), .CI(u5_mult_82_SUMB_9__37_), .CO(
        u5_mult_82_CARRYB_10__36_), .S(u5_mult_82_SUMB_10__36_) );
  FA_X1 u5_mult_82_S2_10_35 ( .A(u5_mult_82_ab_10__35_), .B(
        u5_mult_82_CARRYB_9__35_), .CI(u5_mult_82_SUMB_9__36_), .CO(
        u5_mult_82_CARRYB_10__35_), .S(u5_mult_82_SUMB_10__35_) );
  FA_X1 u5_mult_82_S2_10_34 ( .A(u5_mult_82_ab_10__34_), .B(
        u5_mult_82_CARRYB_9__34_), .CI(u5_mult_82_SUMB_9__35_), .CO(
        u5_mult_82_CARRYB_10__34_), .S(u5_mult_82_SUMB_10__34_) );
  FA_X1 u5_mult_82_S2_10_33 ( .A(u5_mult_82_ab_10__33_), .B(
        u5_mult_82_CARRYB_9__33_), .CI(u5_mult_82_SUMB_9__34_), .CO(
        u5_mult_82_CARRYB_10__33_), .S(u5_mult_82_SUMB_10__33_) );
  FA_X1 u5_mult_82_S2_10_32 ( .A(u5_mult_82_ab_10__32_), .B(
        u5_mult_82_CARRYB_9__32_), .CI(u5_mult_82_SUMB_9__33_), .CO(
        u5_mult_82_CARRYB_10__32_), .S(u5_mult_82_SUMB_10__32_) );
  FA_X1 u5_mult_82_S2_10_31 ( .A(u5_mult_82_ab_10__31_), .B(
        u5_mult_82_CARRYB_9__31_), .CI(u5_mult_82_SUMB_9__32_), .CO(
        u5_mult_82_CARRYB_10__31_), .S(u5_mult_82_SUMB_10__31_) );
  FA_X1 u5_mult_82_S2_10_30 ( .A(u5_mult_82_ab_10__30_), .B(
        u5_mult_82_CARRYB_9__30_), .CI(u5_mult_82_SUMB_9__31_), .CO(
        u5_mult_82_CARRYB_10__30_), .S(u5_mult_82_SUMB_10__30_) );
  FA_X1 u5_mult_82_S2_10_29 ( .A(u5_mult_82_ab_10__29_), .B(
        u5_mult_82_CARRYB_9__29_), .CI(u5_mult_82_SUMB_9__30_), .CO(
        u5_mult_82_CARRYB_10__29_), .S(u5_mult_82_SUMB_10__29_) );
  FA_X1 u5_mult_82_S2_10_28 ( .A(u5_mult_82_ab_10__28_), .B(
        u5_mult_82_CARRYB_9__28_), .CI(u5_mult_82_SUMB_9__29_), .CO(
        u5_mult_82_CARRYB_10__28_), .S(u5_mult_82_SUMB_10__28_) );
  FA_X1 u5_mult_82_S2_10_27 ( .A(u5_mult_82_ab_10__27_), .B(
        u5_mult_82_CARRYB_9__27_), .CI(u5_mult_82_SUMB_9__28_), .CO(
        u5_mult_82_CARRYB_10__27_), .S(u5_mult_82_SUMB_10__27_) );
  FA_X1 u5_mult_82_S2_10_26 ( .A(u5_mult_82_ab_10__26_), .B(
        u5_mult_82_CARRYB_9__26_), .CI(u5_mult_82_SUMB_9__27_), .CO(
        u5_mult_82_CARRYB_10__26_), .S(u5_mult_82_SUMB_10__26_) );
  FA_X1 u5_mult_82_S2_10_25 ( .A(u5_mult_82_ab_10__25_), .B(
        u5_mult_82_CARRYB_9__25_), .CI(u5_mult_82_SUMB_9__26_), .CO(
        u5_mult_82_CARRYB_10__25_), .S(u5_mult_82_SUMB_10__25_) );
  FA_X1 u5_mult_82_S2_10_24 ( .A(u5_mult_82_ab_10__24_), .B(
        u5_mult_82_CARRYB_9__24_), .CI(u5_mult_82_SUMB_9__25_), .CO(
        u5_mult_82_CARRYB_10__24_), .S(u5_mult_82_SUMB_10__24_) );
  FA_X1 u5_mult_82_S2_10_23 ( .A(u5_mult_82_ab_10__23_), .B(
        u5_mult_82_CARRYB_9__23_), .CI(u5_mult_82_SUMB_9__24_), .CO(
        u5_mult_82_CARRYB_10__23_), .S(u5_mult_82_SUMB_10__23_) );
  FA_X1 u5_mult_82_S2_10_22 ( .A(u5_mult_82_ab_10__22_), .B(
        u5_mult_82_CARRYB_9__22_), .CI(u5_mult_82_SUMB_9__23_), .CO(
        u5_mult_82_CARRYB_10__22_), .S(u5_mult_82_SUMB_10__22_) );
  FA_X1 u5_mult_82_S2_10_21 ( .A(u5_mult_82_ab_10__21_), .B(
        u5_mult_82_CARRYB_9__21_), .CI(u5_mult_82_SUMB_9__22_), .CO(
        u5_mult_82_CARRYB_10__21_), .S(u5_mult_82_SUMB_10__21_) );
  FA_X1 u5_mult_82_S2_10_20 ( .A(u5_mult_82_ab_10__20_), .B(
        u5_mult_82_CARRYB_9__20_), .CI(u5_mult_82_SUMB_9__21_), .CO(
        u5_mult_82_CARRYB_10__20_), .S(u5_mult_82_SUMB_10__20_) );
  FA_X1 u5_mult_82_S2_10_19 ( .A(u5_mult_82_ab_10__19_), .B(
        u5_mult_82_CARRYB_9__19_), .CI(u5_mult_82_SUMB_9__20_), .CO(
        u5_mult_82_CARRYB_10__19_), .S(u5_mult_82_SUMB_10__19_) );
  FA_X1 u5_mult_82_S2_10_18 ( .A(u5_mult_82_ab_10__18_), .B(
        u5_mult_82_CARRYB_9__18_), .CI(u5_mult_82_SUMB_9__19_), .CO(
        u5_mult_82_CARRYB_10__18_), .S(u5_mult_82_SUMB_10__18_) );
  FA_X1 u5_mult_82_S2_10_17 ( .A(u5_mult_82_ab_10__17_), .B(
        u5_mult_82_CARRYB_9__17_), .CI(u5_mult_82_SUMB_9__18_), .CO(
        u5_mult_82_CARRYB_10__17_), .S(u5_mult_82_SUMB_10__17_) );
  FA_X1 u5_mult_82_S2_10_16 ( .A(u5_mult_82_ab_10__16_), .B(
        u5_mult_82_CARRYB_9__16_), .CI(u5_mult_82_SUMB_9__17_), .CO(
        u5_mult_82_CARRYB_10__16_), .S(u5_mult_82_SUMB_10__16_) );
  FA_X1 u5_mult_82_S2_10_15 ( .A(u5_mult_82_ab_10__15_), .B(
        u5_mult_82_CARRYB_9__15_), .CI(u5_mult_82_SUMB_9__16_), .CO(
        u5_mult_82_CARRYB_10__15_), .S(u5_mult_82_SUMB_10__15_) );
  FA_X1 u5_mult_82_S2_10_14 ( .A(u5_mult_82_ab_10__14_), .B(
        u5_mult_82_CARRYB_9__14_), .CI(u5_mult_82_SUMB_9__15_), .CO(
        u5_mult_82_CARRYB_10__14_), .S(u5_mult_82_SUMB_10__14_) );
  FA_X1 u5_mult_82_S2_10_13 ( .A(u5_mult_82_ab_10__13_), .B(
        u5_mult_82_CARRYB_9__13_), .CI(u5_mult_82_SUMB_9__14_), .CO(
        u5_mult_82_CARRYB_10__13_), .S(u5_mult_82_SUMB_10__13_) );
  FA_X1 u5_mult_82_S2_10_12 ( .A(u5_mult_82_ab_10__12_), .B(
        u5_mult_82_CARRYB_9__12_), .CI(u5_mult_82_SUMB_9__13_), .CO(
        u5_mult_82_CARRYB_10__12_), .S(u5_mult_82_SUMB_10__12_) );
  FA_X1 u5_mult_82_S2_10_11 ( .A(u5_mult_82_ab_10__11_), .B(
        u5_mult_82_CARRYB_9__11_), .CI(u5_mult_82_SUMB_9__12_), .CO(
        u5_mult_82_CARRYB_10__11_), .S(u5_mult_82_SUMB_10__11_) );
  FA_X1 u5_mult_82_S2_10_10 ( .A(u5_mult_82_ab_10__10_), .B(
        u5_mult_82_CARRYB_9__10_), .CI(u5_mult_82_SUMB_9__11_), .CO(
        u5_mult_82_CARRYB_10__10_), .S(u5_mult_82_SUMB_10__10_) );
  FA_X1 u5_mult_82_S2_10_9 ( .A(u5_mult_82_ab_10__9_), .B(
        u5_mult_82_CARRYB_9__9_), .CI(u5_mult_82_SUMB_9__10_), .CO(
        u5_mult_82_CARRYB_10__9_), .S(u5_mult_82_SUMB_10__9_) );
  FA_X1 u5_mult_82_S2_10_8 ( .A(u5_mult_82_ab_10__8_), .B(
        u5_mult_82_CARRYB_9__8_), .CI(u5_mult_82_SUMB_9__9_), .CO(
        u5_mult_82_CARRYB_10__8_), .S(u5_mult_82_SUMB_10__8_) );
  FA_X1 u5_mult_82_S2_10_7 ( .A(u5_mult_82_ab_10__7_), .B(
        u5_mult_82_CARRYB_9__7_), .CI(u5_mult_82_SUMB_9__8_), .CO(
        u5_mult_82_CARRYB_10__7_), .S(u5_mult_82_SUMB_10__7_) );
  FA_X1 u5_mult_82_S2_10_6 ( .A(u5_mult_82_ab_10__6_), .B(
        u5_mult_82_CARRYB_9__6_), .CI(u5_mult_82_SUMB_9__7_), .CO(
        u5_mult_82_CARRYB_10__6_), .S(u5_mult_82_SUMB_10__6_) );
  FA_X1 u5_mult_82_S2_10_5 ( .A(u5_mult_82_ab_10__5_), .B(
        u5_mult_82_CARRYB_9__5_), .CI(u5_mult_82_SUMB_9__6_), .CO(
        u5_mult_82_CARRYB_10__5_), .S(u5_mult_82_SUMB_10__5_) );
  FA_X1 u5_mult_82_S2_10_4 ( .A(u5_mult_82_ab_10__4_), .B(
        u5_mult_82_CARRYB_9__4_), .CI(u5_mult_82_SUMB_9__5_), .CO(
        u5_mult_82_CARRYB_10__4_), .S(u5_mult_82_SUMB_10__4_) );
  FA_X1 u5_mult_82_S2_10_3 ( .A(u5_mult_82_ab_10__3_), .B(
        u5_mult_82_CARRYB_9__3_), .CI(u5_mult_82_SUMB_9__4_), .CO(
        u5_mult_82_CARRYB_10__3_), .S(u5_mult_82_SUMB_10__3_) );
  FA_X1 u5_mult_82_S2_10_2 ( .A(u5_mult_82_ab_10__2_), .B(
        u5_mult_82_CARRYB_9__2_), .CI(u5_mult_82_SUMB_9__3_), .CO(
        u5_mult_82_CARRYB_10__2_), .S(u5_mult_82_SUMB_10__2_) );
  FA_X1 u5_mult_82_S2_10_1 ( .A(u5_mult_82_ab_10__1_), .B(
        u5_mult_82_CARRYB_9__1_), .CI(u5_mult_82_SUMB_9__2_), .CO(
        u5_mult_82_CARRYB_10__1_), .S(u5_mult_82_SUMB_10__1_) );
  FA_X1 u5_mult_82_S1_10_0 ( .A(u5_mult_82_ab_10__0_), .B(
        u5_mult_82_CARRYB_9__0_), .CI(u5_mult_82_SUMB_9__1_), .CO(
        u5_mult_82_CARRYB_10__0_), .S(u5_N10) );
  FA_X1 u5_mult_82_S3_11_51 ( .A(u5_mult_82_ab_11__51_), .B(
        u5_mult_82_CARRYB_10__51_), .CI(u5_mult_82_ab_10__52_), .CO(
        u5_mult_82_CARRYB_11__51_), .S(u5_mult_82_SUMB_11__51_) );
  FA_X1 u5_mult_82_S2_11_50 ( .A(u5_mult_82_ab_11__50_), .B(
        u5_mult_82_CARRYB_10__50_), .CI(u5_mult_82_SUMB_10__51_), .CO(
        u5_mult_82_CARRYB_11__50_), .S(u5_mult_82_SUMB_11__50_) );
  FA_X1 u5_mult_82_S2_11_49 ( .A(u5_mult_82_ab_11__49_), .B(
        u5_mult_82_CARRYB_10__49_), .CI(u5_mult_82_SUMB_10__50_), .CO(
        u5_mult_82_CARRYB_11__49_), .S(u5_mult_82_SUMB_11__49_) );
  FA_X1 u5_mult_82_S2_11_48 ( .A(u5_mult_82_ab_11__48_), .B(
        u5_mult_82_CARRYB_10__48_), .CI(u5_mult_82_SUMB_10__49_), .CO(
        u5_mult_82_CARRYB_11__48_), .S(u5_mult_82_SUMB_11__48_) );
  FA_X1 u5_mult_82_S2_11_47 ( .A(u5_mult_82_ab_11__47_), .B(
        u5_mult_82_CARRYB_10__47_), .CI(u5_mult_82_SUMB_10__48_), .CO(
        u5_mult_82_CARRYB_11__47_), .S(u5_mult_82_SUMB_11__47_) );
  FA_X1 u5_mult_82_S2_11_46 ( .A(u5_mult_82_ab_11__46_), .B(
        u5_mult_82_CARRYB_10__46_), .CI(u5_mult_82_SUMB_10__47_), .CO(
        u5_mult_82_CARRYB_11__46_), .S(u5_mult_82_SUMB_11__46_) );
  FA_X1 u5_mult_82_S2_11_45 ( .A(u5_mult_82_ab_11__45_), .B(
        u5_mult_82_CARRYB_10__45_), .CI(u5_mult_82_SUMB_10__46_), .CO(
        u5_mult_82_CARRYB_11__45_), .S(u5_mult_82_SUMB_11__45_) );
  FA_X1 u5_mult_82_S2_11_44 ( .A(u5_mult_82_ab_11__44_), .B(
        u5_mult_82_CARRYB_10__44_), .CI(u5_mult_82_SUMB_10__45_), .CO(
        u5_mult_82_CARRYB_11__44_), .S(u5_mult_82_SUMB_11__44_) );
  FA_X1 u5_mult_82_S2_11_43 ( .A(u5_mult_82_ab_11__43_), .B(
        u5_mult_82_CARRYB_10__43_), .CI(u5_mult_82_SUMB_10__44_), .CO(
        u5_mult_82_CARRYB_11__43_), .S(u5_mult_82_SUMB_11__43_) );
  FA_X1 u5_mult_82_S2_11_42 ( .A(u5_mult_82_ab_11__42_), .B(
        u5_mult_82_CARRYB_10__42_), .CI(u5_mult_82_SUMB_10__43_), .CO(
        u5_mult_82_CARRYB_11__42_), .S(u5_mult_82_SUMB_11__42_) );
  FA_X1 u5_mult_82_S2_11_41 ( .A(u5_mult_82_ab_11__41_), .B(
        u5_mult_82_CARRYB_10__41_), .CI(u5_mult_82_SUMB_10__42_), .CO(
        u5_mult_82_CARRYB_11__41_), .S(u5_mult_82_SUMB_11__41_) );
  FA_X1 u5_mult_82_S2_11_40 ( .A(u5_mult_82_ab_11__40_), .B(
        u5_mult_82_CARRYB_10__40_), .CI(u5_mult_82_SUMB_10__41_), .CO(
        u5_mult_82_CARRYB_11__40_), .S(u5_mult_82_SUMB_11__40_) );
  FA_X1 u5_mult_82_S2_11_39 ( .A(u5_mult_82_ab_11__39_), .B(
        u5_mult_82_CARRYB_10__39_), .CI(u5_mult_82_SUMB_10__40_), .CO(
        u5_mult_82_CARRYB_11__39_), .S(u5_mult_82_SUMB_11__39_) );
  FA_X1 u5_mult_82_S2_11_38 ( .A(u5_mult_82_ab_11__38_), .B(
        u5_mult_82_CARRYB_10__38_), .CI(u5_mult_82_SUMB_10__39_), .CO(
        u5_mult_82_CARRYB_11__38_), .S(u5_mult_82_SUMB_11__38_) );
  FA_X1 u5_mult_82_S2_11_37 ( .A(u5_mult_82_ab_11__37_), .B(
        u5_mult_82_CARRYB_10__37_), .CI(u5_mult_82_SUMB_10__38_), .CO(
        u5_mult_82_CARRYB_11__37_), .S(u5_mult_82_SUMB_11__37_) );
  FA_X1 u5_mult_82_S2_11_36 ( .A(u5_mult_82_ab_11__36_), .B(
        u5_mult_82_CARRYB_10__36_), .CI(u5_mult_82_SUMB_10__37_), .CO(
        u5_mult_82_CARRYB_11__36_), .S(u5_mult_82_SUMB_11__36_) );
  FA_X1 u5_mult_82_S2_11_35 ( .A(u5_mult_82_ab_11__35_), .B(
        u5_mult_82_CARRYB_10__35_), .CI(u5_mult_82_SUMB_10__36_), .CO(
        u5_mult_82_CARRYB_11__35_), .S(u5_mult_82_SUMB_11__35_) );
  FA_X1 u5_mult_82_S2_11_34 ( .A(u5_mult_82_ab_11__34_), .B(
        u5_mult_82_CARRYB_10__34_), .CI(u5_mult_82_SUMB_10__35_), .CO(
        u5_mult_82_CARRYB_11__34_), .S(u5_mult_82_SUMB_11__34_) );
  FA_X1 u5_mult_82_S2_11_33 ( .A(u5_mult_82_ab_11__33_), .B(
        u5_mult_82_CARRYB_10__33_), .CI(u5_mult_82_SUMB_10__34_), .CO(
        u5_mult_82_CARRYB_11__33_), .S(u5_mult_82_SUMB_11__33_) );
  FA_X1 u5_mult_82_S2_11_32 ( .A(u5_mult_82_ab_11__32_), .B(
        u5_mult_82_CARRYB_10__32_), .CI(u5_mult_82_SUMB_10__33_), .CO(
        u5_mult_82_CARRYB_11__32_), .S(u5_mult_82_SUMB_11__32_) );
  FA_X1 u5_mult_82_S2_11_31 ( .A(u5_mult_82_ab_11__31_), .B(
        u5_mult_82_CARRYB_10__31_), .CI(u5_mult_82_SUMB_10__32_), .CO(
        u5_mult_82_CARRYB_11__31_), .S(u5_mult_82_SUMB_11__31_) );
  FA_X1 u5_mult_82_S2_11_30 ( .A(u5_mult_82_ab_11__30_), .B(
        u5_mult_82_CARRYB_10__30_), .CI(u5_mult_82_SUMB_10__31_), .CO(
        u5_mult_82_CARRYB_11__30_), .S(u5_mult_82_SUMB_11__30_) );
  FA_X1 u5_mult_82_S2_11_29 ( .A(u5_mult_82_ab_11__29_), .B(
        u5_mult_82_CARRYB_10__29_), .CI(u5_mult_82_SUMB_10__30_), .CO(
        u5_mult_82_CARRYB_11__29_), .S(u5_mult_82_SUMB_11__29_) );
  FA_X1 u5_mult_82_S2_11_28 ( .A(u5_mult_82_ab_11__28_), .B(
        u5_mult_82_CARRYB_10__28_), .CI(u5_mult_82_SUMB_10__29_), .CO(
        u5_mult_82_CARRYB_11__28_), .S(u5_mult_82_SUMB_11__28_) );
  FA_X1 u5_mult_82_S2_11_27 ( .A(u5_mult_82_ab_11__27_), .B(
        u5_mult_82_CARRYB_10__27_), .CI(u5_mult_82_SUMB_10__28_), .CO(
        u5_mult_82_CARRYB_11__27_), .S(u5_mult_82_SUMB_11__27_) );
  FA_X1 u5_mult_82_S2_11_26 ( .A(u5_mult_82_ab_11__26_), .B(
        u5_mult_82_CARRYB_10__26_), .CI(u5_mult_82_SUMB_10__27_), .CO(
        u5_mult_82_CARRYB_11__26_), .S(u5_mult_82_SUMB_11__26_) );
  FA_X1 u5_mult_82_S2_11_25 ( .A(u5_mult_82_ab_11__25_), .B(
        u5_mult_82_CARRYB_10__25_), .CI(u5_mult_82_SUMB_10__26_), .CO(
        u5_mult_82_CARRYB_11__25_), .S(u5_mult_82_SUMB_11__25_) );
  FA_X1 u5_mult_82_S2_11_24 ( .A(u5_mult_82_ab_11__24_), .B(
        u5_mult_82_CARRYB_10__24_), .CI(u5_mult_82_SUMB_10__25_), .CO(
        u5_mult_82_CARRYB_11__24_), .S(u5_mult_82_SUMB_11__24_) );
  FA_X1 u5_mult_82_S2_11_23 ( .A(u5_mult_82_ab_11__23_), .B(
        u5_mult_82_CARRYB_10__23_), .CI(u5_mult_82_SUMB_10__24_), .CO(
        u5_mult_82_CARRYB_11__23_), .S(u5_mult_82_SUMB_11__23_) );
  FA_X1 u5_mult_82_S2_11_22 ( .A(u5_mult_82_ab_11__22_), .B(
        u5_mult_82_CARRYB_10__22_), .CI(u5_mult_82_SUMB_10__23_), .CO(
        u5_mult_82_CARRYB_11__22_), .S(u5_mult_82_SUMB_11__22_) );
  FA_X1 u5_mult_82_S2_11_21 ( .A(u5_mult_82_ab_11__21_), .B(
        u5_mult_82_CARRYB_10__21_), .CI(u5_mult_82_SUMB_10__22_), .CO(
        u5_mult_82_CARRYB_11__21_), .S(u5_mult_82_SUMB_11__21_) );
  FA_X1 u5_mult_82_S2_11_20 ( .A(u5_mult_82_ab_11__20_), .B(
        u5_mult_82_CARRYB_10__20_), .CI(u5_mult_82_SUMB_10__21_), .CO(
        u5_mult_82_CARRYB_11__20_), .S(u5_mult_82_SUMB_11__20_) );
  FA_X1 u5_mult_82_S2_11_19 ( .A(u5_mult_82_ab_11__19_), .B(
        u5_mult_82_CARRYB_10__19_), .CI(u5_mult_82_SUMB_10__20_), .CO(
        u5_mult_82_CARRYB_11__19_), .S(u5_mult_82_SUMB_11__19_) );
  FA_X1 u5_mult_82_S2_11_18 ( .A(u5_mult_82_ab_11__18_), .B(
        u5_mult_82_CARRYB_10__18_), .CI(u5_mult_82_SUMB_10__19_), .CO(
        u5_mult_82_CARRYB_11__18_), .S(u5_mult_82_SUMB_11__18_) );
  FA_X1 u5_mult_82_S2_11_17 ( .A(u5_mult_82_ab_11__17_), .B(
        u5_mult_82_CARRYB_10__17_), .CI(u5_mult_82_SUMB_10__18_), .CO(
        u5_mult_82_CARRYB_11__17_), .S(u5_mult_82_SUMB_11__17_) );
  FA_X1 u5_mult_82_S2_11_16 ( .A(u5_mult_82_ab_11__16_), .B(
        u5_mult_82_CARRYB_10__16_), .CI(u5_mult_82_SUMB_10__17_), .CO(
        u5_mult_82_CARRYB_11__16_), .S(u5_mult_82_SUMB_11__16_) );
  FA_X1 u5_mult_82_S2_11_15 ( .A(u5_mult_82_ab_11__15_), .B(
        u5_mult_82_CARRYB_10__15_), .CI(u5_mult_82_SUMB_10__16_), .CO(
        u5_mult_82_CARRYB_11__15_), .S(u5_mult_82_SUMB_11__15_) );
  FA_X1 u5_mult_82_S2_11_14 ( .A(u5_mult_82_ab_11__14_), .B(
        u5_mult_82_CARRYB_10__14_), .CI(u5_mult_82_SUMB_10__15_), .CO(
        u5_mult_82_CARRYB_11__14_), .S(u5_mult_82_SUMB_11__14_) );
  FA_X1 u5_mult_82_S2_11_13 ( .A(u5_mult_82_ab_11__13_), .B(
        u5_mult_82_CARRYB_10__13_), .CI(u5_mult_82_SUMB_10__14_), .CO(
        u5_mult_82_CARRYB_11__13_), .S(u5_mult_82_SUMB_11__13_) );
  FA_X1 u5_mult_82_S2_11_12 ( .A(u5_mult_82_ab_11__12_), .B(
        u5_mult_82_CARRYB_10__12_), .CI(u5_mult_82_SUMB_10__13_), .CO(
        u5_mult_82_CARRYB_11__12_), .S(u5_mult_82_SUMB_11__12_) );
  FA_X1 u5_mult_82_S2_11_11 ( .A(u5_mult_82_ab_11__11_), .B(
        u5_mult_82_CARRYB_10__11_), .CI(u5_mult_82_SUMB_10__12_), .CO(
        u5_mult_82_CARRYB_11__11_), .S(u5_mult_82_SUMB_11__11_) );
  FA_X1 u5_mult_82_S2_11_10 ( .A(u5_mult_82_ab_11__10_), .B(
        u5_mult_82_CARRYB_10__10_), .CI(u5_mult_82_SUMB_10__11_), .CO(
        u5_mult_82_CARRYB_11__10_), .S(u5_mult_82_SUMB_11__10_) );
  FA_X1 u5_mult_82_S2_11_9 ( .A(u5_mult_82_ab_11__9_), .B(
        u5_mult_82_CARRYB_10__9_), .CI(u5_mult_82_SUMB_10__10_), .CO(
        u5_mult_82_CARRYB_11__9_), .S(u5_mult_82_SUMB_11__9_) );
  FA_X1 u5_mult_82_S2_11_8 ( .A(u5_mult_82_ab_11__8_), .B(
        u5_mult_82_CARRYB_10__8_), .CI(u5_mult_82_SUMB_10__9_), .CO(
        u5_mult_82_CARRYB_11__8_), .S(u5_mult_82_SUMB_11__8_) );
  FA_X1 u5_mult_82_S2_11_7 ( .A(u5_mult_82_ab_11__7_), .B(
        u5_mult_82_CARRYB_10__7_), .CI(u5_mult_82_SUMB_10__8_), .CO(
        u5_mult_82_CARRYB_11__7_), .S(u5_mult_82_SUMB_11__7_) );
  FA_X1 u5_mult_82_S2_11_6 ( .A(u5_mult_82_ab_11__6_), .B(
        u5_mult_82_CARRYB_10__6_), .CI(u5_mult_82_SUMB_10__7_), .CO(
        u5_mult_82_CARRYB_11__6_), .S(u5_mult_82_SUMB_11__6_) );
  FA_X1 u5_mult_82_S2_11_5 ( .A(u5_mult_82_ab_11__5_), .B(
        u5_mult_82_CARRYB_10__5_), .CI(u5_mult_82_SUMB_10__6_), .CO(
        u5_mult_82_CARRYB_11__5_), .S(u5_mult_82_SUMB_11__5_) );
  FA_X1 u5_mult_82_S2_11_4 ( .A(u5_mult_82_ab_11__4_), .B(
        u5_mult_82_CARRYB_10__4_), .CI(u5_mult_82_SUMB_10__5_), .CO(
        u5_mult_82_CARRYB_11__4_), .S(u5_mult_82_SUMB_11__4_) );
  FA_X1 u5_mult_82_S2_11_3 ( .A(u5_mult_82_ab_11__3_), .B(
        u5_mult_82_CARRYB_10__3_), .CI(u5_mult_82_SUMB_10__4_), .CO(
        u5_mult_82_CARRYB_11__3_), .S(u5_mult_82_SUMB_11__3_) );
  FA_X1 u5_mult_82_S2_11_2 ( .A(u5_mult_82_ab_11__2_), .B(
        u5_mult_82_CARRYB_10__2_), .CI(u5_mult_82_SUMB_10__3_), .CO(
        u5_mult_82_CARRYB_11__2_), .S(u5_mult_82_SUMB_11__2_) );
  FA_X1 u5_mult_82_S2_11_1 ( .A(u5_mult_82_ab_11__1_), .B(
        u5_mult_82_CARRYB_10__1_), .CI(u5_mult_82_SUMB_10__2_), .CO(
        u5_mult_82_CARRYB_11__1_), .S(u5_mult_82_SUMB_11__1_) );
  FA_X1 u5_mult_82_S1_11_0 ( .A(u5_mult_82_ab_11__0_), .B(
        u5_mult_82_CARRYB_10__0_), .CI(u5_mult_82_SUMB_10__1_), .CO(
        u5_mult_82_CARRYB_11__0_), .S(u5_N11) );
  FA_X1 u5_mult_82_S3_12_51 ( .A(u5_mult_82_ab_12__51_), .B(
        u5_mult_82_CARRYB_11__51_), .CI(u5_mult_82_ab_11__52_), .CO(
        u5_mult_82_CARRYB_12__51_), .S(u5_mult_82_SUMB_12__51_) );
  FA_X1 u5_mult_82_S2_12_50 ( .A(u5_mult_82_ab_12__50_), .B(
        u5_mult_82_CARRYB_11__50_), .CI(u5_mult_82_SUMB_11__51_), .CO(
        u5_mult_82_CARRYB_12__50_), .S(u5_mult_82_SUMB_12__50_) );
  FA_X1 u5_mult_82_S2_12_49 ( .A(u5_mult_82_ab_12__49_), .B(
        u5_mult_82_CARRYB_11__49_), .CI(u5_mult_82_SUMB_11__50_), .CO(
        u5_mult_82_CARRYB_12__49_), .S(u5_mult_82_SUMB_12__49_) );
  FA_X1 u5_mult_82_S2_12_48 ( .A(u5_mult_82_ab_12__48_), .B(
        u5_mult_82_CARRYB_11__48_), .CI(u5_mult_82_SUMB_11__49_), .CO(
        u5_mult_82_CARRYB_12__48_), .S(u5_mult_82_SUMB_12__48_) );
  FA_X1 u5_mult_82_S2_12_47 ( .A(u5_mult_82_ab_12__47_), .B(
        u5_mult_82_CARRYB_11__47_), .CI(u5_mult_82_SUMB_11__48_), .CO(
        u5_mult_82_CARRYB_12__47_), .S(u5_mult_82_SUMB_12__47_) );
  FA_X1 u5_mult_82_S2_12_46 ( .A(u5_mult_82_ab_12__46_), .B(
        u5_mult_82_CARRYB_11__46_), .CI(u5_mult_82_SUMB_11__47_), .CO(
        u5_mult_82_CARRYB_12__46_), .S(u5_mult_82_SUMB_12__46_) );
  FA_X1 u5_mult_82_S2_12_45 ( .A(u5_mult_82_ab_12__45_), .B(
        u5_mult_82_CARRYB_11__45_), .CI(u5_mult_82_SUMB_11__46_), .CO(
        u5_mult_82_CARRYB_12__45_), .S(u5_mult_82_SUMB_12__45_) );
  FA_X1 u5_mult_82_S2_12_44 ( .A(u5_mult_82_ab_12__44_), .B(
        u5_mult_82_CARRYB_11__44_), .CI(u5_mult_82_SUMB_11__45_), .CO(
        u5_mult_82_CARRYB_12__44_), .S(u5_mult_82_SUMB_12__44_) );
  FA_X1 u5_mult_82_S2_12_43 ( .A(u5_mult_82_ab_12__43_), .B(
        u5_mult_82_CARRYB_11__43_), .CI(u5_mult_82_SUMB_11__44_), .CO(
        u5_mult_82_CARRYB_12__43_), .S(u5_mult_82_SUMB_12__43_) );
  FA_X1 u5_mult_82_S2_12_42 ( .A(u5_mult_82_ab_12__42_), .B(
        u5_mult_82_CARRYB_11__42_), .CI(u5_mult_82_SUMB_11__43_), .CO(
        u5_mult_82_CARRYB_12__42_), .S(u5_mult_82_SUMB_12__42_) );
  FA_X1 u5_mult_82_S2_12_41 ( .A(u5_mult_82_ab_12__41_), .B(
        u5_mult_82_CARRYB_11__41_), .CI(u5_mult_82_SUMB_11__42_), .CO(
        u5_mult_82_CARRYB_12__41_), .S(u5_mult_82_SUMB_12__41_) );
  FA_X1 u5_mult_82_S2_12_40 ( .A(u5_mult_82_ab_12__40_), .B(
        u5_mult_82_CARRYB_11__40_), .CI(u5_mult_82_SUMB_11__41_), .CO(
        u5_mult_82_CARRYB_12__40_), .S(u5_mult_82_SUMB_12__40_) );
  FA_X1 u5_mult_82_S2_12_39 ( .A(u5_mult_82_ab_12__39_), .B(
        u5_mult_82_CARRYB_11__39_), .CI(u5_mult_82_SUMB_11__40_), .CO(
        u5_mult_82_CARRYB_12__39_), .S(u5_mult_82_SUMB_12__39_) );
  FA_X1 u5_mult_82_S2_12_38 ( .A(u5_mult_82_ab_12__38_), .B(
        u5_mult_82_CARRYB_11__38_), .CI(u5_mult_82_SUMB_11__39_), .CO(
        u5_mult_82_CARRYB_12__38_), .S(u5_mult_82_SUMB_12__38_) );
  FA_X1 u5_mult_82_S2_12_37 ( .A(u5_mult_82_ab_12__37_), .B(
        u5_mult_82_CARRYB_11__37_), .CI(u5_mult_82_SUMB_11__38_), .CO(
        u5_mult_82_CARRYB_12__37_), .S(u5_mult_82_SUMB_12__37_) );
  FA_X1 u5_mult_82_S2_12_36 ( .A(u5_mult_82_ab_12__36_), .B(
        u5_mult_82_CARRYB_11__36_), .CI(u5_mult_82_SUMB_11__37_), .CO(
        u5_mult_82_CARRYB_12__36_), .S(u5_mult_82_SUMB_12__36_) );
  FA_X1 u5_mult_82_S2_12_35 ( .A(u5_mult_82_ab_12__35_), .B(
        u5_mult_82_CARRYB_11__35_), .CI(u5_mult_82_SUMB_11__36_), .CO(
        u5_mult_82_CARRYB_12__35_), .S(u5_mult_82_SUMB_12__35_) );
  FA_X1 u5_mult_82_S2_12_34 ( .A(u5_mult_82_ab_12__34_), .B(
        u5_mult_82_CARRYB_11__34_), .CI(u5_mult_82_SUMB_11__35_), .CO(
        u5_mult_82_CARRYB_12__34_), .S(u5_mult_82_SUMB_12__34_) );
  FA_X1 u5_mult_82_S2_12_33 ( .A(u5_mult_82_ab_12__33_), .B(
        u5_mult_82_CARRYB_11__33_), .CI(u5_mult_82_SUMB_11__34_), .CO(
        u5_mult_82_CARRYB_12__33_), .S(u5_mult_82_SUMB_12__33_) );
  FA_X1 u5_mult_82_S2_12_32 ( .A(u5_mult_82_ab_12__32_), .B(
        u5_mult_82_CARRYB_11__32_), .CI(u5_mult_82_SUMB_11__33_), .CO(
        u5_mult_82_CARRYB_12__32_), .S(u5_mult_82_SUMB_12__32_) );
  FA_X1 u5_mult_82_S2_12_31 ( .A(u5_mult_82_ab_12__31_), .B(
        u5_mult_82_CARRYB_11__31_), .CI(u5_mult_82_SUMB_11__32_), .CO(
        u5_mult_82_CARRYB_12__31_), .S(u5_mult_82_SUMB_12__31_) );
  FA_X1 u5_mult_82_S2_12_30 ( .A(u5_mult_82_ab_12__30_), .B(
        u5_mult_82_CARRYB_11__30_), .CI(u5_mult_82_SUMB_11__31_), .CO(
        u5_mult_82_CARRYB_12__30_), .S(u5_mult_82_SUMB_12__30_) );
  FA_X1 u5_mult_82_S2_12_29 ( .A(u5_mult_82_ab_12__29_), .B(
        u5_mult_82_CARRYB_11__29_), .CI(u5_mult_82_SUMB_11__30_), .CO(
        u5_mult_82_CARRYB_12__29_), .S(u5_mult_82_SUMB_12__29_) );
  FA_X1 u5_mult_82_S2_12_28 ( .A(u5_mult_82_ab_12__28_), .B(
        u5_mult_82_CARRYB_11__28_), .CI(u5_mult_82_SUMB_11__29_), .CO(
        u5_mult_82_CARRYB_12__28_), .S(u5_mult_82_SUMB_12__28_) );
  FA_X1 u5_mult_82_S2_12_27 ( .A(u5_mult_82_ab_12__27_), .B(
        u5_mult_82_CARRYB_11__27_), .CI(u5_mult_82_SUMB_11__28_), .CO(
        u5_mult_82_CARRYB_12__27_), .S(u5_mult_82_SUMB_12__27_) );
  FA_X1 u5_mult_82_S2_12_26 ( .A(u5_mult_82_ab_12__26_), .B(
        u5_mult_82_CARRYB_11__26_), .CI(u5_mult_82_SUMB_11__27_), .CO(
        u5_mult_82_CARRYB_12__26_), .S(u5_mult_82_SUMB_12__26_) );
  FA_X1 u5_mult_82_S2_12_25 ( .A(u5_mult_82_ab_12__25_), .B(
        u5_mult_82_CARRYB_11__25_), .CI(u5_mult_82_SUMB_11__26_), .CO(
        u5_mult_82_CARRYB_12__25_), .S(u5_mult_82_SUMB_12__25_) );
  FA_X1 u5_mult_82_S2_12_24 ( .A(u5_mult_82_ab_12__24_), .B(
        u5_mult_82_CARRYB_11__24_), .CI(u5_mult_82_SUMB_11__25_), .CO(
        u5_mult_82_CARRYB_12__24_), .S(u5_mult_82_SUMB_12__24_) );
  FA_X1 u5_mult_82_S2_12_23 ( .A(u5_mult_82_ab_12__23_), .B(
        u5_mult_82_CARRYB_11__23_), .CI(u5_mult_82_SUMB_11__24_), .CO(
        u5_mult_82_CARRYB_12__23_), .S(u5_mult_82_SUMB_12__23_) );
  FA_X1 u5_mult_82_S2_12_22 ( .A(u5_mult_82_ab_12__22_), .B(
        u5_mult_82_CARRYB_11__22_), .CI(u5_mult_82_SUMB_11__23_), .CO(
        u5_mult_82_CARRYB_12__22_), .S(u5_mult_82_SUMB_12__22_) );
  FA_X1 u5_mult_82_S2_12_21 ( .A(u5_mult_82_ab_12__21_), .B(
        u5_mult_82_CARRYB_11__21_), .CI(u5_mult_82_SUMB_11__22_), .CO(
        u5_mult_82_CARRYB_12__21_), .S(u5_mult_82_SUMB_12__21_) );
  FA_X1 u5_mult_82_S2_12_20 ( .A(u5_mult_82_ab_12__20_), .B(
        u5_mult_82_CARRYB_11__20_), .CI(u5_mult_82_SUMB_11__21_), .CO(
        u5_mult_82_CARRYB_12__20_), .S(u5_mult_82_SUMB_12__20_) );
  FA_X1 u5_mult_82_S2_12_19 ( .A(u5_mult_82_ab_12__19_), .B(
        u5_mult_82_CARRYB_11__19_), .CI(u5_mult_82_SUMB_11__20_), .CO(
        u5_mult_82_CARRYB_12__19_), .S(u5_mult_82_SUMB_12__19_) );
  FA_X1 u5_mult_82_S2_12_18 ( .A(u5_mult_82_ab_12__18_), .B(
        u5_mult_82_CARRYB_11__18_), .CI(u5_mult_82_SUMB_11__19_), .CO(
        u5_mult_82_CARRYB_12__18_), .S(u5_mult_82_SUMB_12__18_) );
  FA_X1 u5_mult_82_S2_12_17 ( .A(u5_mult_82_ab_12__17_), .B(
        u5_mult_82_CARRYB_11__17_), .CI(u5_mult_82_SUMB_11__18_), .CO(
        u5_mult_82_CARRYB_12__17_), .S(u5_mult_82_SUMB_12__17_) );
  FA_X1 u5_mult_82_S2_12_16 ( .A(u5_mult_82_ab_12__16_), .B(
        u5_mult_82_CARRYB_11__16_), .CI(u5_mult_82_SUMB_11__17_), .CO(
        u5_mult_82_CARRYB_12__16_), .S(u5_mult_82_SUMB_12__16_) );
  FA_X1 u5_mult_82_S2_12_15 ( .A(u5_mult_82_ab_12__15_), .B(
        u5_mult_82_CARRYB_11__15_), .CI(u5_mult_82_SUMB_11__16_), .CO(
        u5_mult_82_CARRYB_12__15_), .S(u5_mult_82_SUMB_12__15_) );
  FA_X1 u5_mult_82_S2_12_14 ( .A(u5_mult_82_ab_12__14_), .B(
        u5_mult_82_CARRYB_11__14_), .CI(u5_mult_82_SUMB_11__15_), .CO(
        u5_mult_82_CARRYB_12__14_), .S(u5_mult_82_SUMB_12__14_) );
  FA_X1 u5_mult_82_S2_12_13 ( .A(u5_mult_82_ab_12__13_), .B(
        u5_mult_82_CARRYB_11__13_), .CI(u5_mult_82_SUMB_11__14_), .CO(
        u5_mult_82_CARRYB_12__13_), .S(u5_mult_82_SUMB_12__13_) );
  FA_X1 u5_mult_82_S2_12_12 ( .A(u5_mult_82_ab_12__12_), .B(
        u5_mult_82_CARRYB_11__12_), .CI(u5_mult_82_SUMB_11__13_), .CO(
        u5_mult_82_CARRYB_12__12_), .S(u5_mult_82_SUMB_12__12_) );
  FA_X1 u5_mult_82_S2_12_11 ( .A(u5_mult_82_ab_12__11_), .B(
        u5_mult_82_CARRYB_11__11_), .CI(u5_mult_82_SUMB_11__12_), .CO(
        u5_mult_82_CARRYB_12__11_), .S(u5_mult_82_SUMB_12__11_) );
  FA_X1 u5_mult_82_S2_12_10 ( .A(u5_mult_82_ab_12__10_), .B(
        u5_mult_82_CARRYB_11__10_), .CI(u5_mult_82_SUMB_11__11_), .CO(
        u5_mult_82_CARRYB_12__10_), .S(u5_mult_82_SUMB_12__10_) );
  FA_X1 u5_mult_82_S2_12_9 ( .A(u5_mult_82_ab_12__9_), .B(
        u5_mult_82_CARRYB_11__9_), .CI(u5_mult_82_SUMB_11__10_), .CO(
        u5_mult_82_CARRYB_12__9_), .S(u5_mult_82_SUMB_12__9_) );
  FA_X1 u5_mult_82_S2_12_8 ( .A(u5_mult_82_ab_12__8_), .B(
        u5_mult_82_CARRYB_11__8_), .CI(u5_mult_82_SUMB_11__9_), .CO(
        u5_mult_82_CARRYB_12__8_), .S(u5_mult_82_SUMB_12__8_) );
  FA_X1 u5_mult_82_S2_12_7 ( .A(u5_mult_82_ab_12__7_), .B(
        u5_mult_82_CARRYB_11__7_), .CI(u5_mult_82_SUMB_11__8_), .CO(
        u5_mult_82_CARRYB_12__7_), .S(u5_mult_82_SUMB_12__7_) );
  FA_X1 u5_mult_82_S2_12_6 ( .A(u5_mult_82_ab_12__6_), .B(
        u5_mult_82_CARRYB_11__6_), .CI(u5_mult_82_SUMB_11__7_), .CO(
        u5_mult_82_CARRYB_12__6_), .S(u5_mult_82_SUMB_12__6_) );
  FA_X1 u5_mult_82_S2_12_5 ( .A(u5_mult_82_ab_12__5_), .B(
        u5_mult_82_CARRYB_11__5_), .CI(u5_mult_82_SUMB_11__6_), .CO(
        u5_mult_82_CARRYB_12__5_), .S(u5_mult_82_SUMB_12__5_) );
  FA_X1 u5_mult_82_S2_12_4 ( .A(u5_mult_82_ab_12__4_), .B(
        u5_mult_82_CARRYB_11__4_), .CI(u5_mult_82_SUMB_11__5_), .CO(
        u5_mult_82_CARRYB_12__4_), .S(u5_mult_82_SUMB_12__4_) );
  FA_X1 u5_mult_82_S2_12_3 ( .A(u5_mult_82_ab_12__3_), .B(
        u5_mult_82_CARRYB_11__3_), .CI(u5_mult_82_SUMB_11__4_), .CO(
        u5_mult_82_CARRYB_12__3_), .S(u5_mult_82_SUMB_12__3_) );
  FA_X1 u5_mult_82_S2_12_2 ( .A(u5_mult_82_ab_12__2_), .B(
        u5_mult_82_CARRYB_11__2_), .CI(u5_mult_82_SUMB_11__3_), .CO(
        u5_mult_82_CARRYB_12__2_), .S(u5_mult_82_SUMB_12__2_) );
  FA_X1 u5_mult_82_S2_12_1 ( .A(u5_mult_82_ab_12__1_), .B(
        u5_mult_82_CARRYB_11__1_), .CI(u5_mult_82_SUMB_11__2_), .CO(
        u5_mult_82_CARRYB_12__1_), .S(u5_mult_82_SUMB_12__1_) );
  FA_X1 u5_mult_82_S1_12_0 ( .A(u5_mult_82_ab_12__0_), .B(
        u5_mult_82_CARRYB_11__0_), .CI(u5_mult_82_SUMB_11__1_), .CO(
        u5_mult_82_CARRYB_12__0_), .S(u5_N12) );
  FA_X1 u5_mult_82_S3_13_51 ( .A(u5_mult_82_ab_13__51_), .B(
        u5_mult_82_CARRYB_12__51_), .CI(u5_mult_82_ab_12__52_), .CO(
        u5_mult_82_CARRYB_13__51_), .S(u5_mult_82_SUMB_13__51_) );
  FA_X1 u5_mult_82_S2_13_50 ( .A(u5_mult_82_ab_13__50_), .B(
        u5_mult_82_CARRYB_12__50_), .CI(u5_mult_82_SUMB_12__51_), .CO(
        u5_mult_82_CARRYB_13__50_), .S(u5_mult_82_SUMB_13__50_) );
  FA_X1 u5_mult_82_S2_13_49 ( .A(u5_mult_82_ab_13__49_), .B(
        u5_mult_82_CARRYB_12__49_), .CI(u5_mult_82_SUMB_12__50_), .CO(
        u5_mult_82_CARRYB_13__49_), .S(u5_mult_82_SUMB_13__49_) );
  FA_X1 u5_mult_82_S2_13_48 ( .A(u5_mult_82_ab_13__48_), .B(
        u5_mult_82_CARRYB_12__48_), .CI(u5_mult_82_SUMB_12__49_), .CO(
        u5_mult_82_CARRYB_13__48_), .S(u5_mult_82_SUMB_13__48_) );
  FA_X1 u5_mult_82_S2_13_47 ( .A(u5_mult_82_ab_13__47_), .B(
        u5_mult_82_CARRYB_12__47_), .CI(u5_mult_82_SUMB_12__48_), .CO(
        u5_mult_82_CARRYB_13__47_), .S(u5_mult_82_SUMB_13__47_) );
  FA_X1 u5_mult_82_S2_13_46 ( .A(u5_mult_82_ab_13__46_), .B(
        u5_mult_82_CARRYB_12__46_), .CI(u5_mult_82_SUMB_12__47_), .CO(
        u5_mult_82_CARRYB_13__46_), .S(u5_mult_82_SUMB_13__46_) );
  FA_X1 u5_mult_82_S2_13_45 ( .A(u5_mult_82_ab_13__45_), .B(
        u5_mult_82_CARRYB_12__45_), .CI(u5_mult_82_SUMB_12__46_), .CO(
        u5_mult_82_CARRYB_13__45_), .S(u5_mult_82_SUMB_13__45_) );
  FA_X1 u5_mult_82_S2_13_44 ( .A(u5_mult_82_ab_13__44_), .B(
        u5_mult_82_CARRYB_12__44_), .CI(u5_mult_82_SUMB_12__45_), .CO(
        u5_mult_82_CARRYB_13__44_), .S(u5_mult_82_SUMB_13__44_) );
  FA_X1 u5_mult_82_S2_13_43 ( .A(u5_mult_82_ab_13__43_), .B(
        u5_mult_82_CARRYB_12__43_), .CI(u5_mult_82_SUMB_12__44_), .CO(
        u5_mult_82_CARRYB_13__43_), .S(u5_mult_82_SUMB_13__43_) );
  FA_X1 u5_mult_82_S2_13_42 ( .A(u5_mult_82_ab_13__42_), .B(
        u5_mult_82_CARRYB_12__42_), .CI(u5_mult_82_SUMB_12__43_), .CO(
        u5_mult_82_CARRYB_13__42_), .S(u5_mult_82_SUMB_13__42_) );
  FA_X1 u5_mult_82_S2_13_41 ( .A(u5_mult_82_ab_13__41_), .B(
        u5_mult_82_CARRYB_12__41_), .CI(u5_mult_82_SUMB_12__42_), .CO(
        u5_mult_82_CARRYB_13__41_), .S(u5_mult_82_SUMB_13__41_) );
  FA_X1 u5_mult_82_S2_13_40 ( .A(u5_mult_82_ab_13__40_), .B(
        u5_mult_82_CARRYB_12__40_), .CI(u5_mult_82_SUMB_12__41_), .CO(
        u5_mult_82_CARRYB_13__40_), .S(u5_mult_82_SUMB_13__40_) );
  FA_X1 u5_mult_82_S2_13_39 ( .A(u5_mult_82_ab_13__39_), .B(
        u5_mult_82_CARRYB_12__39_), .CI(u5_mult_82_SUMB_12__40_), .CO(
        u5_mult_82_CARRYB_13__39_), .S(u5_mult_82_SUMB_13__39_) );
  FA_X1 u5_mult_82_S2_13_38 ( .A(u5_mult_82_ab_13__38_), .B(
        u5_mult_82_CARRYB_12__38_), .CI(u5_mult_82_SUMB_12__39_), .CO(
        u5_mult_82_CARRYB_13__38_), .S(u5_mult_82_SUMB_13__38_) );
  FA_X1 u5_mult_82_S2_13_37 ( .A(u5_mult_82_ab_13__37_), .B(
        u5_mult_82_CARRYB_12__37_), .CI(u5_mult_82_SUMB_12__38_), .CO(
        u5_mult_82_CARRYB_13__37_), .S(u5_mult_82_SUMB_13__37_) );
  FA_X1 u5_mult_82_S2_13_36 ( .A(u5_mult_82_ab_13__36_), .B(
        u5_mult_82_CARRYB_12__36_), .CI(u5_mult_82_SUMB_12__37_), .CO(
        u5_mult_82_CARRYB_13__36_), .S(u5_mult_82_SUMB_13__36_) );
  FA_X1 u5_mult_82_S2_13_35 ( .A(u5_mult_82_ab_13__35_), .B(
        u5_mult_82_CARRYB_12__35_), .CI(u5_mult_82_SUMB_12__36_), .CO(
        u5_mult_82_CARRYB_13__35_), .S(u5_mult_82_SUMB_13__35_) );
  FA_X1 u5_mult_82_S2_13_34 ( .A(u5_mult_82_ab_13__34_), .B(
        u5_mult_82_CARRYB_12__34_), .CI(u5_mult_82_SUMB_12__35_), .CO(
        u5_mult_82_CARRYB_13__34_), .S(u5_mult_82_SUMB_13__34_) );
  FA_X1 u5_mult_82_S2_13_33 ( .A(u5_mult_82_ab_13__33_), .B(
        u5_mult_82_CARRYB_12__33_), .CI(u5_mult_82_SUMB_12__34_), .CO(
        u5_mult_82_CARRYB_13__33_), .S(u5_mult_82_SUMB_13__33_) );
  FA_X1 u5_mult_82_S2_13_32 ( .A(u5_mult_82_ab_13__32_), .B(
        u5_mult_82_CARRYB_12__32_), .CI(u5_mult_82_SUMB_12__33_), .CO(
        u5_mult_82_CARRYB_13__32_), .S(u5_mult_82_SUMB_13__32_) );
  FA_X1 u5_mult_82_S2_13_31 ( .A(u5_mult_82_ab_13__31_), .B(
        u5_mult_82_CARRYB_12__31_), .CI(u5_mult_82_SUMB_12__32_), .CO(
        u5_mult_82_CARRYB_13__31_), .S(u5_mult_82_SUMB_13__31_) );
  FA_X1 u5_mult_82_S2_13_30 ( .A(u5_mult_82_ab_13__30_), .B(
        u5_mult_82_CARRYB_12__30_), .CI(u5_mult_82_SUMB_12__31_), .CO(
        u5_mult_82_CARRYB_13__30_), .S(u5_mult_82_SUMB_13__30_) );
  FA_X1 u5_mult_82_S2_13_29 ( .A(u5_mult_82_ab_13__29_), .B(
        u5_mult_82_CARRYB_12__29_), .CI(u5_mult_82_SUMB_12__30_), .CO(
        u5_mult_82_CARRYB_13__29_), .S(u5_mult_82_SUMB_13__29_) );
  FA_X1 u5_mult_82_S2_13_28 ( .A(u5_mult_82_ab_13__28_), .B(
        u5_mult_82_CARRYB_12__28_), .CI(u5_mult_82_SUMB_12__29_), .CO(
        u5_mult_82_CARRYB_13__28_), .S(u5_mult_82_SUMB_13__28_) );
  FA_X1 u5_mult_82_S2_13_27 ( .A(u5_mult_82_ab_13__27_), .B(
        u5_mult_82_CARRYB_12__27_), .CI(u5_mult_82_SUMB_12__28_), .CO(
        u5_mult_82_CARRYB_13__27_), .S(u5_mult_82_SUMB_13__27_) );
  FA_X1 u5_mult_82_S2_13_26 ( .A(u5_mult_82_ab_13__26_), .B(
        u5_mult_82_CARRYB_12__26_), .CI(u5_mult_82_SUMB_12__27_), .CO(
        u5_mult_82_CARRYB_13__26_), .S(u5_mult_82_SUMB_13__26_) );
  FA_X1 u5_mult_82_S2_13_25 ( .A(u5_mult_82_ab_13__25_), .B(
        u5_mult_82_CARRYB_12__25_), .CI(u5_mult_82_SUMB_12__26_), .CO(
        u5_mult_82_CARRYB_13__25_), .S(u5_mult_82_SUMB_13__25_) );
  FA_X1 u5_mult_82_S2_13_24 ( .A(u5_mult_82_ab_13__24_), .B(
        u5_mult_82_CARRYB_12__24_), .CI(u5_mult_82_SUMB_12__25_), .CO(
        u5_mult_82_CARRYB_13__24_), .S(u5_mult_82_SUMB_13__24_) );
  FA_X1 u5_mult_82_S2_13_23 ( .A(u5_mult_82_ab_13__23_), .B(
        u5_mult_82_CARRYB_12__23_), .CI(u5_mult_82_SUMB_12__24_), .CO(
        u5_mult_82_CARRYB_13__23_), .S(u5_mult_82_SUMB_13__23_) );
  FA_X1 u5_mult_82_S2_13_22 ( .A(u5_mult_82_ab_13__22_), .B(
        u5_mult_82_CARRYB_12__22_), .CI(u5_mult_82_SUMB_12__23_), .CO(
        u5_mult_82_CARRYB_13__22_), .S(u5_mult_82_SUMB_13__22_) );
  FA_X1 u5_mult_82_S2_13_21 ( .A(u5_mult_82_ab_13__21_), .B(
        u5_mult_82_CARRYB_12__21_), .CI(u5_mult_82_SUMB_12__22_), .CO(
        u5_mult_82_CARRYB_13__21_), .S(u5_mult_82_SUMB_13__21_) );
  FA_X1 u5_mult_82_S2_13_20 ( .A(u5_mult_82_ab_13__20_), .B(
        u5_mult_82_CARRYB_12__20_), .CI(u5_mult_82_SUMB_12__21_), .CO(
        u5_mult_82_CARRYB_13__20_), .S(u5_mult_82_SUMB_13__20_) );
  FA_X1 u5_mult_82_S2_13_19 ( .A(u5_mult_82_ab_13__19_), .B(
        u5_mult_82_CARRYB_12__19_), .CI(u5_mult_82_SUMB_12__20_), .CO(
        u5_mult_82_CARRYB_13__19_), .S(u5_mult_82_SUMB_13__19_) );
  FA_X1 u5_mult_82_S2_13_18 ( .A(u5_mult_82_ab_13__18_), .B(
        u5_mult_82_CARRYB_12__18_), .CI(u5_mult_82_SUMB_12__19_), .CO(
        u5_mult_82_CARRYB_13__18_), .S(u5_mult_82_SUMB_13__18_) );
  FA_X1 u5_mult_82_S2_13_17 ( .A(u5_mult_82_ab_13__17_), .B(
        u5_mult_82_CARRYB_12__17_), .CI(u5_mult_82_SUMB_12__18_), .CO(
        u5_mult_82_CARRYB_13__17_), .S(u5_mult_82_SUMB_13__17_) );
  FA_X1 u5_mult_82_S2_13_16 ( .A(u5_mult_82_ab_13__16_), .B(
        u5_mult_82_CARRYB_12__16_), .CI(u5_mult_82_SUMB_12__17_), .CO(
        u5_mult_82_CARRYB_13__16_), .S(u5_mult_82_SUMB_13__16_) );
  FA_X1 u5_mult_82_S2_13_15 ( .A(u5_mult_82_ab_13__15_), .B(
        u5_mult_82_CARRYB_12__15_), .CI(u5_mult_82_SUMB_12__16_), .CO(
        u5_mult_82_CARRYB_13__15_), .S(u5_mult_82_SUMB_13__15_) );
  FA_X1 u5_mult_82_S2_13_14 ( .A(u5_mult_82_ab_13__14_), .B(
        u5_mult_82_CARRYB_12__14_), .CI(u5_mult_82_SUMB_12__15_), .CO(
        u5_mult_82_CARRYB_13__14_), .S(u5_mult_82_SUMB_13__14_) );
  FA_X1 u5_mult_82_S2_13_13 ( .A(u5_mult_82_ab_13__13_), .B(
        u5_mult_82_CARRYB_12__13_), .CI(u5_mult_82_SUMB_12__14_), .CO(
        u5_mult_82_CARRYB_13__13_), .S(u5_mult_82_SUMB_13__13_) );
  FA_X1 u5_mult_82_S2_13_12 ( .A(u5_mult_82_ab_13__12_), .B(
        u5_mult_82_CARRYB_12__12_), .CI(u5_mult_82_SUMB_12__13_), .CO(
        u5_mult_82_CARRYB_13__12_), .S(u5_mult_82_SUMB_13__12_) );
  FA_X1 u5_mult_82_S2_13_11 ( .A(u5_mult_82_ab_13__11_), .B(
        u5_mult_82_CARRYB_12__11_), .CI(u5_mult_82_SUMB_12__12_), .CO(
        u5_mult_82_CARRYB_13__11_), .S(u5_mult_82_SUMB_13__11_) );
  FA_X1 u5_mult_82_S2_13_10 ( .A(u5_mult_82_ab_13__10_), .B(
        u5_mult_82_CARRYB_12__10_), .CI(u5_mult_82_SUMB_12__11_), .CO(
        u5_mult_82_CARRYB_13__10_), .S(u5_mult_82_SUMB_13__10_) );
  FA_X1 u5_mult_82_S2_13_9 ( .A(u5_mult_82_ab_13__9_), .B(
        u5_mult_82_CARRYB_12__9_), .CI(u5_mult_82_SUMB_12__10_), .CO(
        u5_mult_82_CARRYB_13__9_), .S(u5_mult_82_SUMB_13__9_) );
  FA_X1 u5_mult_82_S2_13_8 ( .A(u5_mult_82_ab_13__8_), .B(
        u5_mult_82_CARRYB_12__8_), .CI(u5_mult_82_SUMB_12__9_), .CO(
        u5_mult_82_CARRYB_13__8_), .S(u5_mult_82_SUMB_13__8_) );
  FA_X1 u5_mult_82_S2_13_7 ( .A(u5_mult_82_ab_13__7_), .B(
        u5_mult_82_CARRYB_12__7_), .CI(u5_mult_82_SUMB_12__8_), .CO(
        u5_mult_82_CARRYB_13__7_), .S(u5_mult_82_SUMB_13__7_) );
  FA_X1 u5_mult_82_S2_13_6 ( .A(u5_mult_82_ab_13__6_), .B(
        u5_mult_82_CARRYB_12__6_), .CI(u5_mult_82_SUMB_12__7_), .CO(
        u5_mult_82_CARRYB_13__6_), .S(u5_mult_82_SUMB_13__6_) );
  FA_X1 u5_mult_82_S2_13_5 ( .A(u5_mult_82_ab_13__5_), .B(
        u5_mult_82_CARRYB_12__5_), .CI(u5_mult_82_SUMB_12__6_), .CO(
        u5_mult_82_CARRYB_13__5_), .S(u5_mult_82_SUMB_13__5_) );
  FA_X1 u5_mult_82_S2_13_4 ( .A(u5_mult_82_ab_13__4_), .B(
        u5_mult_82_CARRYB_12__4_), .CI(u5_mult_82_SUMB_12__5_), .CO(
        u5_mult_82_CARRYB_13__4_), .S(u5_mult_82_SUMB_13__4_) );
  FA_X1 u5_mult_82_S2_13_3 ( .A(u5_mult_82_ab_13__3_), .B(
        u5_mult_82_CARRYB_12__3_), .CI(u5_mult_82_SUMB_12__4_), .CO(
        u5_mult_82_CARRYB_13__3_), .S(u5_mult_82_SUMB_13__3_) );
  FA_X1 u5_mult_82_S2_13_2 ( .A(u5_mult_82_ab_13__2_), .B(
        u5_mult_82_CARRYB_12__2_), .CI(u5_mult_82_SUMB_12__3_), .CO(
        u5_mult_82_CARRYB_13__2_), .S(u5_mult_82_SUMB_13__2_) );
  FA_X1 u5_mult_82_S2_13_1 ( .A(u5_mult_82_ab_13__1_), .B(
        u5_mult_82_CARRYB_12__1_), .CI(u5_mult_82_SUMB_12__2_), .CO(
        u5_mult_82_CARRYB_13__1_), .S(u5_mult_82_SUMB_13__1_) );
  FA_X1 u5_mult_82_S1_13_0 ( .A(u5_mult_82_ab_13__0_), .B(
        u5_mult_82_CARRYB_12__0_), .CI(u5_mult_82_SUMB_12__1_), .CO(
        u5_mult_82_CARRYB_13__0_), .S(u5_N13) );
  FA_X1 u5_mult_82_S3_14_51 ( .A(u5_mult_82_ab_14__51_), .B(
        u5_mult_82_CARRYB_13__51_), .CI(u5_mult_82_ab_13__52_), .CO(
        u5_mult_82_CARRYB_14__51_), .S(u5_mult_82_SUMB_14__51_) );
  FA_X1 u5_mult_82_S2_14_50 ( .A(u5_mult_82_ab_14__50_), .B(
        u5_mult_82_CARRYB_13__50_), .CI(u5_mult_82_SUMB_13__51_), .CO(
        u5_mult_82_CARRYB_14__50_), .S(u5_mult_82_SUMB_14__50_) );
  FA_X1 u5_mult_82_S2_14_49 ( .A(u5_mult_82_ab_14__49_), .B(
        u5_mult_82_CARRYB_13__49_), .CI(u5_mult_82_SUMB_13__50_), .CO(
        u5_mult_82_CARRYB_14__49_), .S(u5_mult_82_SUMB_14__49_) );
  FA_X1 u5_mult_82_S2_14_48 ( .A(u5_mult_82_ab_14__48_), .B(
        u5_mult_82_CARRYB_13__48_), .CI(u5_mult_82_SUMB_13__49_), .CO(
        u5_mult_82_CARRYB_14__48_), .S(u5_mult_82_SUMB_14__48_) );
  FA_X1 u5_mult_82_S2_14_47 ( .A(u5_mult_82_ab_14__47_), .B(
        u5_mult_82_CARRYB_13__47_), .CI(u5_mult_82_SUMB_13__48_), .CO(
        u5_mult_82_CARRYB_14__47_), .S(u5_mult_82_SUMB_14__47_) );
  FA_X1 u5_mult_82_S2_14_46 ( .A(u5_mult_82_ab_14__46_), .B(
        u5_mult_82_CARRYB_13__46_), .CI(u5_mult_82_SUMB_13__47_), .CO(
        u5_mult_82_CARRYB_14__46_), .S(u5_mult_82_SUMB_14__46_) );
  FA_X1 u5_mult_82_S2_14_45 ( .A(u5_mult_82_ab_14__45_), .B(
        u5_mult_82_CARRYB_13__45_), .CI(u5_mult_82_SUMB_13__46_), .CO(
        u5_mult_82_CARRYB_14__45_), .S(u5_mult_82_SUMB_14__45_) );
  FA_X1 u5_mult_82_S2_14_44 ( .A(u5_mult_82_ab_14__44_), .B(
        u5_mult_82_CARRYB_13__44_), .CI(u5_mult_82_SUMB_13__45_), .CO(
        u5_mult_82_CARRYB_14__44_), .S(u5_mult_82_SUMB_14__44_) );
  FA_X1 u5_mult_82_S2_14_43 ( .A(u5_mult_82_ab_14__43_), .B(
        u5_mult_82_CARRYB_13__43_), .CI(u5_mult_82_SUMB_13__44_), .CO(
        u5_mult_82_CARRYB_14__43_), .S(u5_mult_82_SUMB_14__43_) );
  FA_X1 u5_mult_82_S2_14_42 ( .A(u5_mult_82_ab_14__42_), .B(
        u5_mult_82_CARRYB_13__42_), .CI(u5_mult_82_SUMB_13__43_), .CO(
        u5_mult_82_CARRYB_14__42_), .S(u5_mult_82_SUMB_14__42_) );
  FA_X1 u5_mult_82_S2_14_41 ( .A(u5_mult_82_ab_14__41_), .B(
        u5_mult_82_CARRYB_13__41_), .CI(u5_mult_82_SUMB_13__42_), .CO(
        u5_mult_82_CARRYB_14__41_), .S(u5_mult_82_SUMB_14__41_) );
  FA_X1 u5_mult_82_S2_14_40 ( .A(u5_mult_82_ab_14__40_), .B(
        u5_mult_82_CARRYB_13__40_), .CI(u5_mult_82_SUMB_13__41_), .CO(
        u5_mult_82_CARRYB_14__40_), .S(u5_mult_82_SUMB_14__40_) );
  FA_X1 u5_mult_82_S2_14_39 ( .A(u5_mult_82_ab_14__39_), .B(
        u5_mult_82_CARRYB_13__39_), .CI(u5_mult_82_SUMB_13__40_), .CO(
        u5_mult_82_CARRYB_14__39_), .S(u5_mult_82_SUMB_14__39_) );
  FA_X1 u5_mult_82_S2_14_38 ( .A(u5_mult_82_ab_14__38_), .B(
        u5_mult_82_CARRYB_13__38_), .CI(u5_mult_82_SUMB_13__39_), .CO(
        u5_mult_82_CARRYB_14__38_), .S(u5_mult_82_SUMB_14__38_) );
  FA_X1 u5_mult_82_S2_14_37 ( .A(u5_mult_82_ab_14__37_), .B(
        u5_mult_82_CARRYB_13__37_), .CI(u5_mult_82_SUMB_13__38_), .CO(
        u5_mult_82_CARRYB_14__37_), .S(u5_mult_82_SUMB_14__37_) );
  FA_X1 u5_mult_82_S2_14_36 ( .A(u5_mult_82_ab_14__36_), .B(
        u5_mult_82_CARRYB_13__36_), .CI(u5_mult_82_SUMB_13__37_), .CO(
        u5_mult_82_CARRYB_14__36_), .S(u5_mult_82_SUMB_14__36_) );
  FA_X1 u5_mult_82_S2_14_35 ( .A(u5_mult_82_ab_14__35_), .B(
        u5_mult_82_CARRYB_13__35_), .CI(u5_mult_82_SUMB_13__36_), .CO(
        u5_mult_82_CARRYB_14__35_), .S(u5_mult_82_SUMB_14__35_) );
  FA_X1 u5_mult_82_S2_14_34 ( .A(u5_mult_82_ab_14__34_), .B(
        u5_mult_82_CARRYB_13__34_), .CI(u5_mult_82_SUMB_13__35_), .CO(
        u5_mult_82_CARRYB_14__34_), .S(u5_mult_82_SUMB_14__34_) );
  FA_X1 u5_mult_82_S2_14_33 ( .A(u5_mult_82_ab_14__33_), .B(
        u5_mult_82_CARRYB_13__33_), .CI(u5_mult_82_SUMB_13__34_), .CO(
        u5_mult_82_CARRYB_14__33_), .S(u5_mult_82_SUMB_14__33_) );
  FA_X1 u5_mult_82_S2_14_32 ( .A(u5_mult_82_ab_14__32_), .B(
        u5_mult_82_CARRYB_13__32_), .CI(u5_mult_82_SUMB_13__33_), .CO(
        u5_mult_82_CARRYB_14__32_), .S(u5_mult_82_SUMB_14__32_) );
  FA_X1 u5_mult_82_S2_14_31 ( .A(u5_mult_82_ab_14__31_), .B(
        u5_mult_82_CARRYB_13__31_), .CI(u5_mult_82_SUMB_13__32_), .CO(
        u5_mult_82_CARRYB_14__31_), .S(u5_mult_82_SUMB_14__31_) );
  FA_X1 u5_mult_82_S2_14_30 ( .A(u5_mult_82_ab_14__30_), .B(
        u5_mult_82_CARRYB_13__30_), .CI(u5_mult_82_SUMB_13__31_), .CO(
        u5_mult_82_CARRYB_14__30_), .S(u5_mult_82_SUMB_14__30_) );
  FA_X1 u5_mult_82_S2_14_29 ( .A(u5_mult_82_ab_14__29_), .B(
        u5_mult_82_CARRYB_13__29_), .CI(u5_mult_82_SUMB_13__30_), .CO(
        u5_mult_82_CARRYB_14__29_), .S(u5_mult_82_SUMB_14__29_) );
  FA_X1 u5_mult_82_S2_14_28 ( .A(u5_mult_82_ab_14__28_), .B(
        u5_mult_82_CARRYB_13__28_), .CI(u5_mult_82_SUMB_13__29_), .CO(
        u5_mult_82_CARRYB_14__28_), .S(u5_mult_82_SUMB_14__28_) );
  FA_X1 u5_mult_82_S2_14_27 ( .A(u5_mult_82_ab_14__27_), .B(
        u5_mult_82_CARRYB_13__27_), .CI(u5_mult_82_SUMB_13__28_), .CO(
        u5_mult_82_CARRYB_14__27_), .S(u5_mult_82_SUMB_14__27_) );
  FA_X1 u5_mult_82_S2_14_26 ( .A(u5_mult_82_ab_14__26_), .B(
        u5_mult_82_CARRYB_13__26_), .CI(u5_mult_82_SUMB_13__27_), .CO(
        u5_mult_82_CARRYB_14__26_), .S(u5_mult_82_SUMB_14__26_) );
  FA_X1 u5_mult_82_S2_14_25 ( .A(u5_mult_82_ab_14__25_), .B(
        u5_mult_82_CARRYB_13__25_), .CI(u5_mult_82_SUMB_13__26_), .CO(
        u5_mult_82_CARRYB_14__25_), .S(u5_mult_82_SUMB_14__25_) );
  FA_X1 u5_mult_82_S2_14_24 ( .A(u5_mult_82_ab_14__24_), .B(
        u5_mult_82_CARRYB_13__24_), .CI(u5_mult_82_SUMB_13__25_), .CO(
        u5_mult_82_CARRYB_14__24_), .S(u5_mult_82_SUMB_14__24_) );
  FA_X1 u5_mult_82_S2_14_23 ( .A(u5_mult_82_ab_14__23_), .B(
        u5_mult_82_CARRYB_13__23_), .CI(u5_mult_82_SUMB_13__24_), .CO(
        u5_mult_82_CARRYB_14__23_), .S(u5_mult_82_SUMB_14__23_) );
  FA_X1 u5_mult_82_S2_14_22 ( .A(u5_mult_82_ab_14__22_), .B(
        u5_mult_82_CARRYB_13__22_), .CI(u5_mult_82_SUMB_13__23_), .CO(
        u5_mult_82_CARRYB_14__22_), .S(u5_mult_82_SUMB_14__22_) );
  FA_X1 u5_mult_82_S2_14_21 ( .A(u5_mult_82_ab_14__21_), .B(
        u5_mult_82_CARRYB_13__21_), .CI(u5_mult_82_SUMB_13__22_), .CO(
        u5_mult_82_CARRYB_14__21_), .S(u5_mult_82_SUMB_14__21_) );
  FA_X1 u5_mult_82_S2_14_20 ( .A(u5_mult_82_ab_14__20_), .B(
        u5_mult_82_CARRYB_13__20_), .CI(u5_mult_82_SUMB_13__21_), .CO(
        u5_mult_82_CARRYB_14__20_), .S(u5_mult_82_SUMB_14__20_) );
  FA_X1 u5_mult_82_S2_14_19 ( .A(u5_mult_82_ab_14__19_), .B(
        u5_mult_82_CARRYB_13__19_), .CI(u5_mult_82_SUMB_13__20_), .CO(
        u5_mult_82_CARRYB_14__19_), .S(u5_mult_82_SUMB_14__19_) );
  FA_X1 u5_mult_82_S2_14_18 ( .A(u5_mult_82_ab_14__18_), .B(
        u5_mult_82_CARRYB_13__18_), .CI(u5_mult_82_SUMB_13__19_), .CO(
        u5_mult_82_CARRYB_14__18_), .S(u5_mult_82_SUMB_14__18_) );
  FA_X1 u5_mult_82_S2_14_17 ( .A(u5_mult_82_ab_14__17_), .B(
        u5_mult_82_CARRYB_13__17_), .CI(u5_mult_82_SUMB_13__18_), .CO(
        u5_mult_82_CARRYB_14__17_), .S(u5_mult_82_SUMB_14__17_) );
  FA_X1 u5_mult_82_S2_14_16 ( .A(u5_mult_82_ab_14__16_), .B(
        u5_mult_82_CARRYB_13__16_), .CI(u5_mult_82_SUMB_13__17_), .CO(
        u5_mult_82_CARRYB_14__16_), .S(u5_mult_82_SUMB_14__16_) );
  FA_X1 u5_mult_82_S2_14_15 ( .A(u5_mult_82_ab_14__15_), .B(
        u5_mult_82_CARRYB_13__15_), .CI(u5_mult_82_SUMB_13__16_), .CO(
        u5_mult_82_CARRYB_14__15_), .S(u5_mult_82_SUMB_14__15_) );
  FA_X1 u5_mult_82_S2_14_14 ( .A(u5_mult_82_ab_14__14_), .B(
        u5_mult_82_CARRYB_13__14_), .CI(u5_mult_82_SUMB_13__15_), .CO(
        u5_mult_82_CARRYB_14__14_), .S(u5_mult_82_SUMB_14__14_) );
  FA_X1 u5_mult_82_S2_14_13 ( .A(u5_mult_82_ab_14__13_), .B(
        u5_mult_82_CARRYB_13__13_), .CI(u5_mult_82_SUMB_13__14_), .CO(
        u5_mult_82_CARRYB_14__13_), .S(u5_mult_82_SUMB_14__13_) );
  FA_X1 u5_mult_82_S2_14_12 ( .A(u5_mult_82_ab_14__12_), .B(
        u5_mult_82_CARRYB_13__12_), .CI(u5_mult_82_SUMB_13__13_), .CO(
        u5_mult_82_CARRYB_14__12_), .S(u5_mult_82_SUMB_14__12_) );
  FA_X1 u5_mult_82_S2_14_11 ( .A(u5_mult_82_ab_14__11_), .B(
        u5_mult_82_CARRYB_13__11_), .CI(u5_mult_82_SUMB_13__12_), .CO(
        u5_mult_82_CARRYB_14__11_), .S(u5_mult_82_SUMB_14__11_) );
  FA_X1 u5_mult_82_S2_14_10 ( .A(u5_mult_82_ab_14__10_), .B(
        u5_mult_82_CARRYB_13__10_), .CI(u5_mult_82_SUMB_13__11_), .CO(
        u5_mult_82_CARRYB_14__10_), .S(u5_mult_82_SUMB_14__10_) );
  FA_X1 u5_mult_82_S2_14_9 ( .A(u5_mult_82_ab_14__9_), .B(
        u5_mult_82_CARRYB_13__9_), .CI(u5_mult_82_SUMB_13__10_), .CO(
        u5_mult_82_CARRYB_14__9_), .S(u5_mult_82_SUMB_14__9_) );
  FA_X1 u5_mult_82_S2_14_8 ( .A(u5_mult_82_ab_14__8_), .B(
        u5_mult_82_CARRYB_13__8_), .CI(u5_mult_82_SUMB_13__9_), .CO(
        u5_mult_82_CARRYB_14__8_), .S(u5_mult_82_SUMB_14__8_) );
  FA_X1 u5_mult_82_S2_14_7 ( .A(u5_mult_82_ab_14__7_), .B(
        u5_mult_82_CARRYB_13__7_), .CI(u5_mult_82_SUMB_13__8_), .CO(
        u5_mult_82_CARRYB_14__7_), .S(u5_mult_82_SUMB_14__7_) );
  FA_X1 u5_mult_82_S2_14_6 ( .A(u5_mult_82_ab_14__6_), .B(
        u5_mult_82_CARRYB_13__6_), .CI(u5_mult_82_SUMB_13__7_), .CO(
        u5_mult_82_CARRYB_14__6_), .S(u5_mult_82_SUMB_14__6_) );
  FA_X1 u5_mult_82_S2_14_5 ( .A(u5_mult_82_ab_14__5_), .B(
        u5_mult_82_CARRYB_13__5_), .CI(u5_mult_82_SUMB_13__6_), .CO(
        u5_mult_82_CARRYB_14__5_), .S(u5_mult_82_SUMB_14__5_) );
  FA_X1 u5_mult_82_S2_14_4 ( .A(u5_mult_82_ab_14__4_), .B(
        u5_mult_82_CARRYB_13__4_), .CI(u5_mult_82_SUMB_13__5_), .CO(
        u5_mult_82_CARRYB_14__4_), .S(u5_mult_82_SUMB_14__4_) );
  FA_X1 u5_mult_82_S2_14_3 ( .A(u5_mult_82_ab_14__3_), .B(
        u5_mult_82_CARRYB_13__3_), .CI(u5_mult_82_SUMB_13__4_), .CO(
        u5_mult_82_CARRYB_14__3_), .S(u5_mult_82_SUMB_14__3_) );
  FA_X1 u5_mult_82_S2_14_2 ( .A(u5_mult_82_ab_14__2_), .B(
        u5_mult_82_CARRYB_13__2_), .CI(u5_mult_82_SUMB_13__3_), .CO(
        u5_mult_82_CARRYB_14__2_), .S(u5_mult_82_SUMB_14__2_) );
  FA_X1 u5_mult_82_S2_14_1 ( .A(u5_mult_82_ab_14__1_), .B(
        u5_mult_82_CARRYB_13__1_), .CI(u5_mult_82_SUMB_13__2_), .CO(
        u5_mult_82_CARRYB_14__1_), .S(u5_mult_82_SUMB_14__1_) );
  FA_X1 u5_mult_82_S1_14_0 ( .A(u5_mult_82_ab_14__0_), .B(
        u5_mult_82_CARRYB_13__0_), .CI(u5_mult_82_SUMB_13__1_), .CO(
        u5_mult_82_CARRYB_14__0_), .S(u5_N14) );
  FA_X1 u5_mult_82_S3_15_51 ( .A(u5_mult_82_ab_15__51_), .B(
        u5_mult_82_CARRYB_14__51_), .CI(u5_mult_82_ab_14__52_), .CO(
        u5_mult_82_CARRYB_15__51_), .S(u5_mult_82_SUMB_15__51_) );
  FA_X1 u5_mult_82_S2_15_50 ( .A(u5_mult_82_ab_15__50_), .B(
        u5_mult_82_CARRYB_14__50_), .CI(u5_mult_82_SUMB_14__51_), .CO(
        u5_mult_82_CARRYB_15__50_), .S(u5_mult_82_SUMB_15__50_) );
  FA_X1 u5_mult_82_S2_15_49 ( .A(u5_mult_82_ab_15__49_), .B(
        u5_mult_82_CARRYB_14__49_), .CI(u5_mult_82_SUMB_14__50_), .CO(
        u5_mult_82_CARRYB_15__49_), .S(u5_mult_82_SUMB_15__49_) );
  FA_X1 u5_mult_82_S2_15_48 ( .A(u5_mult_82_ab_15__48_), .B(
        u5_mult_82_CARRYB_14__48_), .CI(u5_mult_82_SUMB_14__49_), .CO(
        u5_mult_82_CARRYB_15__48_), .S(u5_mult_82_SUMB_15__48_) );
  FA_X1 u5_mult_82_S2_15_47 ( .A(u5_mult_82_ab_15__47_), .B(
        u5_mult_82_CARRYB_14__47_), .CI(u5_mult_82_SUMB_14__48_), .CO(
        u5_mult_82_CARRYB_15__47_), .S(u5_mult_82_SUMB_15__47_) );
  FA_X1 u5_mult_82_S2_15_46 ( .A(u5_mult_82_ab_15__46_), .B(
        u5_mult_82_CARRYB_14__46_), .CI(u5_mult_82_SUMB_14__47_), .CO(
        u5_mult_82_CARRYB_15__46_), .S(u5_mult_82_SUMB_15__46_) );
  FA_X1 u5_mult_82_S2_15_45 ( .A(u5_mult_82_ab_15__45_), .B(
        u5_mult_82_CARRYB_14__45_), .CI(u5_mult_82_SUMB_14__46_), .CO(
        u5_mult_82_CARRYB_15__45_), .S(u5_mult_82_SUMB_15__45_) );
  FA_X1 u5_mult_82_S2_15_44 ( .A(u5_mult_82_ab_15__44_), .B(
        u5_mult_82_CARRYB_14__44_), .CI(u5_mult_82_SUMB_14__45_), .CO(
        u5_mult_82_CARRYB_15__44_), .S(u5_mult_82_SUMB_15__44_) );
  FA_X1 u5_mult_82_S2_15_43 ( .A(u5_mult_82_ab_15__43_), .B(
        u5_mult_82_CARRYB_14__43_), .CI(u5_mult_82_SUMB_14__44_), .CO(
        u5_mult_82_CARRYB_15__43_), .S(u5_mult_82_SUMB_15__43_) );
  FA_X1 u5_mult_82_S2_15_42 ( .A(u5_mult_82_ab_15__42_), .B(
        u5_mult_82_CARRYB_14__42_), .CI(u5_mult_82_SUMB_14__43_), .CO(
        u5_mult_82_CARRYB_15__42_), .S(u5_mult_82_SUMB_15__42_) );
  FA_X1 u5_mult_82_S2_15_41 ( .A(u5_mult_82_ab_15__41_), .B(
        u5_mult_82_CARRYB_14__41_), .CI(u5_mult_82_SUMB_14__42_), .CO(
        u5_mult_82_CARRYB_15__41_), .S(u5_mult_82_SUMB_15__41_) );
  FA_X1 u5_mult_82_S2_15_40 ( .A(u5_mult_82_ab_15__40_), .B(
        u5_mult_82_CARRYB_14__40_), .CI(u5_mult_82_SUMB_14__41_), .CO(
        u5_mult_82_CARRYB_15__40_), .S(u5_mult_82_SUMB_15__40_) );
  FA_X1 u5_mult_82_S2_15_39 ( .A(u5_mult_82_ab_15__39_), .B(
        u5_mult_82_CARRYB_14__39_), .CI(u5_mult_82_SUMB_14__40_), .CO(
        u5_mult_82_CARRYB_15__39_), .S(u5_mult_82_SUMB_15__39_) );
  FA_X1 u5_mult_82_S2_15_38 ( .A(u5_mult_82_ab_15__38_), .B(
        u5_mult_82_CARRYB_14__38_), .CI(u5_mult_82_SUMB_14__39_), .CO(
        u5_mult_82_CARRYB_15__38_), .S(u5_mult_82_SUMB_15__38_) );
  FA_X1 u5_mult_82_S2_15_37 ( .A(u5_mult_82_ab_15__37_), .B(
        u5_mult_82_CARRYB_14__37_), .CI(u5_mult_82_SUMB_14__38_), .CO(
        u5_mult_82_CARRYB_15__37_), .S(u5_mult_82_SUMB_15__37_) );
  FA_X1 u5_mult_82_S2_15_36 ( .A(u5_mult_82_ab_15__36_), .B(
        u5_mult_82_CARRYB_14__36_), .CI(u5_mult_82_SUMB_14__37_), .CO(
        u5_mult_82_CARRYB_15__36_), .S(u5_mult_82_SUMB_15__36_) );
  FA_X1 u5_mult_82_S2_15_35 ( .A(u5_mult_82_ab_15__35_), .B(
        u5_mult_82_CARRYB_14__35_), .CI(u5_mult_82_SUMB_14__36_), .CO(
        u5_mult_82_CARRYB_15__35_), .S(u5_mult_82_SUMB_15__35_) );
  FA_X1 u5_mult_82_S2_15_34 ( .A(u5_mult_82_ab_15__34_), .B(
        u5_mult_82_CARRYB_14__34_), .CI(u5_mult_82_SUMB_14__35_), .CO(
        u5_mult_82_CARRYB_15__34_), .S(u5_mult_82_SUMB_15__34_) );
  FA_X1 u5_mult_82_S2_15_33 ( .A(u5_mult_82_ab_15__33_), .B(
        u5_mult_82_CARRYB_14__33_), .CI(u5_mult_82_SUMB_14__34_), .CO(
        u5_mult_82_CARRYB_15__33_), .S(u5_mult_82_SUMB_15__33_) );
  FA_X1 u5_mult_82_S2_15_32 ( .A(u5_mult_82_ab_15__32_), .B(
        u5_mult_82_CARRYB_14__32_), .CI(u5_mult_82_SUMB_14__33_), .CO(
        u5_mult_82_CARRYB_15__32_), .S(u5_mult_82_SUMB_15__32_) );
  FA_X1 u5_mult_82_S2_15_31 ( .A(u5_mult_82_ab_15__31_), .B(
        u5_mult_82_CARRYB_14__31_), .CI(u5_mult_82_SUMB_14__32_), .CO(
        u5_mult_82_CARRYB_15__31_), .S(u5_mult_82_SUMB_15__31_) );
  FA_X1 u5_mult_82_S2_15_30 ( .A(u5_mult_82_ab_15__30_), .B(
        u5_mult_82_CARRYB_14__30_), .CI(u5_mult_82_SUMB_14__31_), .CO(
        u5_mult_82_CARRYB_15__30_), .S(u5_mult_82_SUMB_15__30_) );
  FA_X1 u5_mult_82_S2_15_29 ( .A(u5_mult_82_ab_15__29_), .B(
        u5_mult_82_CARRYB_14__29_), .CI(u5_mult_82_SUMB_14__30_), .CO(
        u5_mult_82_CARRYB_15__29_), .S(u5_mult_82_SUMB_15__29_) );
  FA_X1 u5_mult_82_S2_15_28 ( .A(u5_mult_82_ab_15__28_), .B(
        u5_mult_82_CARRYB_14__28_), .CI(u5_mult_82_SUMB_14__29_), .CO(
        u5_mult_82_CARRYB_15__28_), .S(u5_mult_82_SUMB_15__28_) );
  FA_X1 u5_mult_82_S2_15_27 ( .A(u5_mult_82_ab_15__27_), .B(
        u5_mult_82_CARRYB_14__27_), .CI(u5_mult_82_SUMB_14__28_), .CO(
        u5_mult_82_CARRYB_15__27_), .S(u5_mult_82_SUMB_15__27_) );
  FA_X1 u5_mult_82_S2_15_26 ( .A(u5_mult_82_ab_15__26_), .B(
        u5_mult_82_CARRYB_14__26_), .CI(u5_mult_82_SUMB_14__27_), .CO(
        u5_mult_82_CARRYB_15__26_), .S(u5_mult_82_SUMB_15__26_) );
  FA_X1 u5_mult_82_S2_15_25 ( .A(u5_mult_82_ab_15__25_), .B(
        u5_mult_82_CARRYB_14__25_), .CI(u5_mult_82_SUMB_14__26_), .CO(
        u5_mult_82_CARRYB_15__25_), .S(u5_mult_82_SUMB_15__25_) );
  FA_X1 u5_mult_82_S2_15_24 ( .A(u5_mult_82_ab_15__24_), .B(
        u5_mult_82_CARRYB_14__24_), .CI(u5_mult_82_SUMB_14__25_), .CO(
        u5_mult_82_CARRYB_15__24_), .S(u5_mult_82_SUMB_15__24_) );
  FA_X1 u5_mult_82_S2_15_23 ( .A(u5_mult_82_ab_15__23_), .B(
        u5_mult_82_CARRYB_14__23_), .CI(u5_mult_82_SUMB_14__24_), .CO(
        u5_mult_82_CARRYB_15__23_), .S(u5_mult_82_SUMB_15__23_) );
  FA_X1 u5_mult_82_S2_15_22 ( .A(u5_mult_82_ab_15__22_), .B(
        u5_mult_82_CARRYB_14__22_), .CI(u5_mult_82_SUMB_14__23_), .CO(
        u5_mult_82_CARRYB_15__22_), .S(u5_mult_82_SUMB_15__22_) );
  FA_X1 u5_mult_82_S2_15_21 ( .A(u5_mult_82_ab_15__21_), .B(
        u5_mult_82_CARRYB_14__21_), .CI(u5_mult_82_SUMB_14__22_), .CO(
        u5_mult_82_CARRYB_15__21_), .S(u5_mult_82_SUMB_15__21_) );
  FA_X1 u5_mult_82_S2_15_20 ( .A(u5_mult_82_ab_15__20_), .B(
        u5_mult_82_CARRYB_14__20_), .CI(u5_mult_82_SUMB_14__21_), .CO(
        u5_mult_82_CARRYB_15__20_), .S(u5_mult_82_SUMB_15__20_) );
  FA_X1 u5_mult_82_S2_15_19 ( .A(u5_mult_82_ab_15__19_), .B(
        u5_mult_82_CARRYB_14__19_), .CI(u5_mult_82_SUMB_14__20_), .CO(
        u5_mult_82_CARRYB_15__19_), .S(u5_mult_82_SUMB_15__19_) );
  FA_X1 u5_mult_82_S2_15_18 ( .A(u5_mult_82_ab_15__18_), .B(
        u5_mult_82_CARRYB_14__18_), .CI(u5_mult_82_SUMB_14__19_), .CO(
        u5_mult_82_CARRYB_15__18_), .S(u5_mult_82_SUMB_15__18_) );
  FA_X1 u5_mult_82_S2_15_17 ( .A(u5_mult_82_ab_15__17_), .B(
        u5_mult_82_CARRYB_14__17_), .CI(u5_mult_82_SUMB_14__18_), .CO(
        u5_mult_82_CARRYB_15__17_), .S(u5_mult_82_SUMB_15__17_) );
  FA_X1 u5_mult_82_S2_15_16 ( .A(u5_mult_82_ab_15__16_), .B(
        u5_mult_82_CARRYB_14__16_), .CI(u5_mult_82_SUMB_14__17_), .CO(
        u5_mult_82_CARRYB_15__16_), .S(u5_mult_82_SUMB_15__16_) );
  FA_X1 u5_mult_82_S2_15_15 ( .A(u5_mult_82_ab_15__15_), .B(
        u5_mult_82_CARRYB_14__15_), .CI(u5_mult_82_SUMB_14__16_), .CO(
        u5_mult_82_CARRYB_15__15_), .S(u5_mult_82_SUMB_15__15_) );
  FA_X1 u5_mult_82_S2_15_14 ( .A(u5_mult_82_ab_15__14_), .B(
        u5_mult_82_CARRYB_14__14_), .CI(u5_mult_82_SUMB_14__15_), .CO(
        u5_mult_82_CARRYB_15__14_), .S(u5_mult_82_SUMB_15__14_) );
  FA_X1 u5_mult_82_S2_15_13 ( .A(u5_mult_82_ab_15__13_), .B(
        u5_mult_82_CARRYB_14__13_), .CI(u5_mult_82_SUMB_14__14_), .CO(
        u5_mult_82_CARRYB_15__13_), .S(u5_mult_82_SUMB_15__13_) );
  FA_X1 u5_mult_82_S2_15_12 ( .A(u5_mult_82_ab_15__12_), .B(
        u5_mult_82_CARRYB_14__12_), .CI(u5_mult_82_SUMB_14__13_), .CO(
        u5_mult_82_CARRYB_15__12_), .S(u5_mult_82_SUMB_15__12_) );
  FA_X1 u5_mult_82_S2_15_11 ( .A(u5_mult_82_ab_15__11_), .B(
        u5_mult_82_CARRYB_14__11_), .CI(u5_mult_82_SUMB_14__12_), .CO(
        u5_mult_82_CARRYB_15__11_), .S(u5_mult_82_SUMB_15__11_) );
  FA_X1 u5_mult_82_S2_15_10 ( .A(u5_mult_82_ab_15__10_), .B(
        u5_mult_82_CARRYB_14__10_), .CI(u5_mult_82_SUMB_14__11_), .CO(
        u5_mult_82_CARRYB_15__10_), .S(u5_mult_82_SUMB_15__10_) );
  FA_X1 u5_mult_82_S2_15_9 ( .A(u5_mult_82_ab_15__9_), .B(
        u5_mult_82_CARRYB_14__9_), .CI(u5_mult_82_SUMB_14__10_), .CO(
        u5_mult_82_CARRYB_15__9_), .S(u5_mult_82_SUMB_15__9_) );
  FA_X1 u5_mult_82_S2_15_8 ( .A(u5_mult_82_ab_15__8_), .B(
        u5_mult_82_CARRYB_14__8_), .CI(u5_mult_82_SUMB_14__9_), .CO(
        u5_mult_82_CARRYB_15__8_), .S(u5_mult_82_SUMB_15__8_) );
  FA_X1 u5_mult_82_S2_15_7 ( .A(u5_mult_82_ab_15__7_), .B(
        u5_mult_82_CARRYB_14__7_), .CI(u5_mult_82_SUMB_14__8_), .CO(
        u5_mult_82_CARRYB_15__7_), .S(u5_mult_82_SUMB_15__7_) );
  FA_X1 u5_mult_82_S2_15_6 ( .A(u5_mult_82_ab_15__6_), .B(
        u5_mult_82_CARRYB_14__6_), .CI(u5_mult_82_SUMB_14__7_), .CO(
        u5_mult_82_CARRYB_15__6_), .S(u5_mult_82_SUMB_15__6_) );
  FA_X1 u5_mult_82_S2_15_5 ( .A(u5_mult_82_ab_15__5_), .B(
        u5_mult_82_CARRYB_14__5_), .CI(u5_mult_82_SUMB_14__6_), .CO(
        u5_mult_82_CARRYB_15__5_), .S(u5_mult_82_SUMB_15__5_) );
  FA_X1 u5_mult_82_S2_15_4 ( .A(u5_mult_82_ab_15__4_), .B(
        u5_mult_82_CARRYB_14__4_), .CI(u5_mult_82_SUMB_14__5_), .CO(
        u5_mult_82_CARRYB_15__4_), .S(u5_mult_82_SUMB_15__4_) );
  FA_X1 u5_mult_82_S2_15_3 ( .A(u5_mult_82_ab_15__3_), .B(
        u5_mult_82_CARRYB_14__3_), .CI(u5_mult_82_SUMB_14__4_), .CO(
        u5_mult_82_CARRYB_15__3_), .S(u5_mult_82_SUMB_15__3_) );
  FA_X1 u5_mult_82_S2_15_2 ( .A(u5_mult_82_ab_15__2_), .B(
        u5_mult_82_CARRYB_14__2_), .CI(u5_mult_82_SUMB_14__3_), .CO(
        u5_mult_82_CARRYB_15__2_), .S(u5_mult_82_SUMB_15__2_) );
  FA_X1 u5_mult_82_S2_15_1 ( .A(u5_mult_82_ab_15__1_), .B(
        u5_mult_82_CARRYB_14__1_), .CI(u5_mult_82_SUMB_14__2_), .CO(
        u5_mult_82_CARRYB_15__1_), .S(u5_mult_82_SUMB_15__1_) );
  FA_X1 u5_mult_82_S1_15_0 ( .A(u5_mult_82_ab_15__0_), .B(
        u5_mult_82_CARRYB_14__0_), .CI(u5_mult_82_SUMB_14__1_), .CO(
        u5_mult_82_CARRYB_15__0_), .S(u5_N15) );
  FA_X1 u5_mult_82_S3_16_51 ( .A(u5_mult_82_ab_16__51_), .B(
        u5_mult_82_CARRYB_15__51_), .CI(u5_mult_82_ab_15__52_), .CO(
        u5_mult_82_CARRYB_16__51_), .S(u5_mult_82_SUMB_16__51_) );
  FA_X1 u5_mult_82_S2_16_50 ( .A(u5_mult_82_ab_16__50_), .B(
        u5_mult_82_CARRYB_15__50_), .CI(u5_mult_82_SUMB_15__51_), .CO(
        u5_mult_82_CARRYB_16__50_), .S(u5_mult_82_SUMB_16__50_) );
  FA_X1 u5_mult_82_S2_16_49 ( .A(u5_mult_82_ab_16__49_), .B(
        u5_mult_82_CARRYB_15__49_), .CI(u5_mult_82_SUMB_15__50_), .CO(
        u5_mult_82_CARRYB_16__49_), .S(u5_mult_82_SUMB_16__49_) );
  FA_X1 u5_mult_82_S2_16_48 ( .A(u5_mult_82_ab_16__48_), .B(
        u5_mult_82_CARRYB_15__48_), .CI(u5_mult_82_SUMB_15__49_), .CO(
        u5_mult_82_CARRYB_16__48_), .S(u5_mult_82_SUMB_16__48_) );
  FA_X1 u5_mult_82_S2_16_47 ( .A(u5_mult_82_ab_16__47_), .B(
        u5_mult_82_CARRYB_15__47_), .CI(u5_mult_82_SUMB_15__48_), .CO(
        u5_mult_82_CARRYB_16__47_), .S(u5_mult_82_SUMB_16__47_) );
  FA_X1 u5_mult_82_S2_16_46 ( .A(u5_mult_82_ab_16__46_), .B(
        u5_mult_82_CARRYB_15__46_), .CI(u5_mult_82_SUMB_15__47_), .CO(
        u5_mult_82_CARRYB_16__46_), .S(u5_mult_82_SUMB_16__46_) );
  FA_X1 u5_mult_82_S2_16_45 ( .A(u5_mult_82_ab_16__45_), .B(
        u5_mult_82_CARRYB_15__45_), .CI(u5_mult_82_SUMB_15__46_), .CO(
        u5_mult_82_CARRYB_16__45_), .S(u5_mult_82_SUMB_16__45_) );
  FA_X1 u5_mult_82_S2_16_44 ( .A(u5_mult_82_ab_16__44_), .B(
        u5_mult_82_CARRYB_15__44_), .CI(u5_mult_82_SUMB_15__45_), .CO(
        u5_mult_82_CARRYB_16__44_), .S(u5_mult_82_SUMB_16__44_) );
  FA_X1 u5_mult_82_S2_16_43 ( .A(u5_mult_82_ab_16__43_), .B(
        u5_mult_82_CARRYB_15__43_), .CI(u5_mult_82_SUMB_15__44_), .CO(
        u5_mult_82_CARRYB_16__43_), .S(u5_mult_82_SUMB_16__43_) );
  FA_X1 u5_mult_82_S2_16_42 ( .A(u5_mult_82_ab_16__42_), .B(
        u5_mult_82_CARRYB_15__42_), .CI(u5_mult_82_SUMB_15__43_), .CO(
        u5_mult_82_CARRYB_16__42_), .S(u5_mult_82_SUMB_16__42_) );
  FA_X1 u5_mult_82_S2_16_41 ( .A(u5_mult_82_ab_16__41_), .B(
        u5_mult_82_CARRYB_15__41_), .CI(u5_mult_82_SUMB_15__42_), .CO(
        u5_mult_82_CARRYB_16__41_), .S(u5_mult_82_SUMB_16__41_) );
  FA_X1 u5_mult_82_S2_16_40 ( .A(u5_mult_82_ab_16__40_), .B(
        u5_mult_82_CARRYB_15__40_), .CI(u5_mult_82_SUMB_15__41_), .CO(
        u5_mult_82_CARRYB_16__40_), .S(u5_mult_82_SUMB_16__40_) );
  FA_X1 u5_mult_82_S2_16_39 ( .A(u5_mult_82_ab_16__39_), .B(
        u5_mult_82_CARRYB_15__39_), .CI(u5_mult_82_SUMB_15__40_), .CO(
        u5_mult_82_CARRYB_16__39_), .S(u5_mult_82_SUMB_16__39_) );
  FA_X1 u5_mult_82_S2_16_38 ( .A(u5_mult_82_ab_16__38_), .B(
        u5_mult_82_CARRYB_15__38_), .CI(u5_mult_82_SUMB_15__39_), .CO(
        u5_mult_82_CARRYB_16__38_), .S(u5_mult_82_SUMB_16__38_) );
  FA_X1 u5_mult_82_S2_16_37 ( .A(u5_mult_82_ab_16__37_), .B(
        u5_mult_82_CARRYB_15__37_), .CI(u5_mult_82_SUMB_15__38_), .CO(
        u5_mult_82_CARRYB_16__37_), .S(u5_mult_82_SUMB_16__37_) );
  FA_X1 u5_mult_82_S2_16_36 ( .A(u5_mult_82_ab_16__36_), .B(
        u5_mult_82_CARRYB_15__36_), .CI(u5_mult_82_SUMB_15__37_), .CO(
        u5_mult_82_CARRYB_16__36_), .S(u5_mult_82_SUMB_16__36_) );
  FA_X1 u5_mult_82_S2_16_35 ( .A(u5_mult_82_ab_16__35_), .B(
        u5_mult_82_CARRYB_15__35_), .CI(u5_mult_82_SUMB_15__36_), .CO(
        u5_mult_82_CARRYB_16__35_), .S(u5_mult_82_SUMB_16__35_) );
  FA_X1 u5_mult_82_S2_16_34 ( .A(u5_mult_82_ab_16__34_), .B(
        u5_mult_82_CARRYB_15__34_), .CI(u5_mult_82_SUMB_15__35_), .CO(
        u5_mult_82_CARRYB_16__34_), .S(u5_mult_82_SUMB_16__34_) );
  FA_X1 u5_mult_82_S2_16_33 ( .A(u5_mult_82_ab_16__33_), .B(
        u5_mult_82_CARRYB_15__33_), .CI(u5_mult_82_SUMB_15__34_), .CO(
        u5_mult_82_CARRYB_16__33_), .S(u5_mult_82_SUMB_16__33_) );
  FA_X1 u5_mult_82_S2_16_32 ( .A(u5_mult_82_ab_16__32_), .B(
        u5_mult_82_CARRYB_15__32_), .CI(u5_mult_82_SUMB_15__33_), .CO(
        u5_mult_82_CARRYB_16__32_), .S(u5_mult_82_SUMB_16__32_) );
  FA_X1 u5_mult_82_S2_16_31 ( .A(u5_mult_82_ab_16__31_), .B(
        u5_mult_82_CARRYB_15__31_), .CI(u5_mult_82_SUMB_15__32_), .CO(
        u5_mult_82_CARRYB_16__31_), .S(u5_mult_82_SUMB_16__31_) );
  FA_X1 u5_mult_82_S2_16_30 ( .A(u5_mult_82_ab_16__30_), .B(
        u5_mult_82_CARRYB_15__30_), .CI(u5_mult_82_SUMB_15__31_), .CO(
        u5_mult_82_CARRYB_16__30_), .S(u5_mult_82_SUMB_16__30_) );
  FA_X1 u5_mult_82_S2_16_29 ( .A(u5_mult_82_ab_16__29_), .B(
        u5_mult_82_CARRYB_15__29_), .CI(u5_mult_82_SUMB_15__30_), .CO(
        u5_mult_82_CARRYB_16__29_), .S(u5_mult_82_SUMB_16__29_) );
  FA_X1 u5_mult_82_S2_16_28 ( .A(u5_mult_82_ab_16__28_), .B(
        u5_mult_82_CARRYB_15__28_), .CI(u5_mult_82_SUMB_15__29_), .CO(
        u5_mult_82_CARRYB_16__28_), .S(u5_mult_82_SUMB_16__28_) );
  FA_X1 u5_mult_82_S2_16_27 ( .A(u5_mult_82_ab_16__27_), .B(
        u5_mult_82_CARRYB_15__27_), .CI(u5_mult_82_SUMB_15__28_), .CO(
        u5_mult_82_CARRYB_16__27_), .S(u5_mult_82_SUMB_16__27_) );
  FA_X1 u5_mult_82_S2_16_26 ( .A(u5_mult_82_ab_16__26_), .B(
        u5_mult_82_CARRYB_15__26_), .CI(u5_mult_82_SUMB_15__27_), .CO(
        u5_mult_82_CARRYB_16__26_), .S(u5_mult_82_SUMB_16__26_) );
  FA_X1 u5_mult_82_S2_16_25 ( .A(u5_mult_82_ab_16__25_), .B(
        u5_mult_82_CARRYB_15__25_), .CI(u5_mult_82_SUMB_15__26_), .CO(
        u5_mult_82_CARRYB_16__25_), .S(u5_mult_82_SUMB_16__25_) );
  FA_X1 u5_mult_82_S2_16_24 ( .A(u5_mult_82_ab_16__24_), .B(
        u5_mult_82_CARRYB_15__24_), .CI(u5_mult_82_SUMB_15__25_), .CO(
        u5_mult_82_CARRYB_16__24_), .S(u5_mult_82_SUMB_16__24_) );
  FA_X1 u5_mult_82_S2_16_23 ( .A(u5_mult_82_ab_16__23_), .B(
        u5_mult_82_CARRYB_15__23_), .CI(u5_mult_82_SUMB_15__24_), .CO(
        u5_mult_82_CARRYB_16__23_), .S(u5_mult_82_SUMB_16__23_) );
  FA_X1 u5_mult_82_S2_16_22 ( .A(u5_mult_82_ab_16__22_), .B(
        u5_mult_82_CARRYB_15__22_), .CI(u5_mult_82_SUMB_15__23_), .CO(
        u5_mult_82_CARRYB_16__22_), .S(u5_mult_82_SUMB_16__22_) );
  FA_X1 u5_mult_82_S2_16_21 ( .A(u5_mult_82_ab_16__21_), .B(
        u5_mult_82_CARRYB_15__21_), .CI(u5_mult_82_SUMB_15__22_), .CO(
        u5_mult_82_CARRYB_16__21_), .S(u5_mult_82_SUMB_16__21_) );
  FA_X1 u5_mult_82_S2_16_20 ( .A(u5_mult_82_ab_16__20_), .B(
        u5_mult_82_CARRYB_15__20_), .CI(u5_mult_82_SUMB_15__21_), .CO(
        u5_mult_82_CARRYB_16__20_), .S(u5_mult_82_SUMB_16__20_) );
  FA_X1 u5_mult_82_S2_16_19 ( .A(u5_mult_82_ab_16__19_), .B(
        u5_mult_82_CARRYB_15__19_), .CI(u5_mult_82_SUMB_15__20_), .CO(
        u5_mult_82_CARRYB_16__19_), .S(u5_mult_82_SUMB_16__19_) );
  FA_X1 u5_mult_82_S2_16_18 ( .A(u5_mult_82_ab_16__18_), .B(
        u5_mult_82_CARRYB_15__18_), .CI(u5_mult_82_SUMB_15__19_), .CO(
        u5_mult_82_CARRYB_16__18_), .S(u5_mult_82_SUMB_16__18_) );
  FA_X1 u5_mult_82_S2_16_17 ( .A(u5_mult_82_ab_16__17_), .B(
        u5_mult_82_CARRYB_15__17_), .CI(u5_mult_82_SUMB_15__18_), .CO(
        u5_mult_82_CARRYB_16__17_), .S(u5_mult_82_SUMB_16__17_) );
  FA_X1 u5_mult_82_S2_16_16 ( .A(u5_mult_82_ab_16__16_), .B(
        u5_mult_82_CARRYB_15__16_), .CI(u5_mult_82_SUMB_15__17_), .CO(
        u5_mult_82_CARRYB_16__16_), .S(u5_mult_82_SUMB_16__16_) );
  FA_X1 u5_mult_82_S2_16_15 ( .A(u5_mult_82_ab_16__15_), .B(
        u5_mult_82_CARRYB_15__15_), .CI(u5_mult_82_SUMB_15__16_), .CO(
        u5_mult_82_CARRYB_16__15_), .S(u5_mult_82_SUMB_16__15_) );
  FA_X1 u5_mult_82_S2_16_14 ( .A(u5_mult_82_ab_16__14_), .B(
        u5_mult_82_CARRYB_15__14_), .CI(u5_mult_82_SUMB_15__15_), .CO(
        u5_mult_82_CARRYB_16__14_), .S(u5_mult_82_SUMB_16__14_) );
  FA_X1 u5_mult_82_S2_16_13 ( .A(u5_mult_82_ab_16__13_), .B(
        u5_mult_82_CARRYB_15__13_), .CI(u5_mult_82_SUMB_15__14_), .CO(
        u5_mult_82_CARRYB_16__13_), .S(u5_mult_82_SUMB_16__13_) );
  FA_X1 u5_mult_82_S2_16_12 ( .A(u5_mult_82_ab_16__12_), .B(
        u5_mult_82_CARRYB_15__12_), .CI(u5_mult_82_SUMB_15__13_), .CO(
        u5_mult_82_CARRYB_16__12_), .S(u5_mult_82_SUMB_16__12_) );
  FA_X1 u5_mult_82_S2_16_11 ( .A(u5_mult_82_ab_16__11_), .B(
        u5_mult_82_CARRYB_15__11_), .CI(u5_mult_82_SUMB_15__12_), .CO(
        u5_mult_82_CARRYB_16__11_), .S(u5_mult_82_SUMB_16__11_) );
  FA_X1 u5_mult_82_S2_16_10 ( .A(u5_mult_82_ab_16__10_), .B(
        u5_mult_82_CARRYB_15__10_), .CI(u5_mult_82_SUMB_15__11_), .CO(
        u5_mult_82_CARRYB_16__10_), .S(u5_mult_82_SUMB_16__10_) );
  FA_X1 u5_mult_82_S2_16_9 ( .A(u5_mult_82_ab_16__9_), .B(
        u5_mult_82_CARRYB_15__9_), .CI(u5_mult_82_SUMB_15__10_), .CO(
        u5_mult_82_CARRYB_16__9_), .S(u5_mult_82_SUMB_16__9_) );
  FA_X1 u5_mult_82_S2_16_8 ( .A(u5_mult_82_ab_16__8_), .B(
        u5_mult_82_CARRYB_15__8_), .CI(u5_mult_82_SUMB_15__9_), .CO(
        u5_mult_82_CARRYB_16__8_), .S(u5_mult_82_SUMB_16__8_) );
  FA_X1 u5_mult_82_S2_16_7 ( .A(u5_mult_82_ab_16__7_), .B(
        u5_mult_82_CARRYB_15__7_), .CI(u5_mult_82_SUMB_15__8_), .CO(
        u5_mult_82_CARRYB_16__7_), .S(u5_mult_82_SUMB_16__7_) );
  FA_X1 u5_mult_82_S2_16_6 ( .A(u5_mult_82_ab_16__6_), .B(
        u5_mult_82_CARRYB_15__6_), .CI(u5_mult_82_SUMB_15__7_), .CO(
        u5_mult_82_CARRYB_16__6_), .S(u5_mult_82_SUMB_16__6_) );
  FA_X1 u5_mult_82_S2_16_5 ( .A(u5_mult_82_ab_16__5_), .B(
        u5_mult_82_CARRYB_15__5_), .CI(u5_mult_82_SUMB_15__6_), .CO(
        u5_mult_82_CARRYB_16__5_), .S(u5_mult_82_SUMB_16__5_) );
  FA_X1 u5_mult_82_S2_16_4 ( .A(u5_mult_82_ab_16__4_), .B(
        u5_mult_82_CARRYB_15__4_), .CI(u5_mult_82_SUMB_15__5_), .CO(
        u5_mult_82_CARRYB_16__4_), .S(u5_mult_82_SUMB_16__4_) );
  FA_X1 u5_mult_82_S2_16_3 ( .A(u5_mult_82_ab_16__3_), .B(
        u5_mult_82_CARRYB_15__3_), .CI(u5_mult_82_SUMB_15__4_), .CO(
        u5_mult_82_CARRYB_16__3_), .S(u5_mult_82_SUMB_16__3_) );
  FA_X1 u5_mult_82_S2_16_2 ( .A(u5_mult_82_ab_16__2_), .B(
        u5_mult_82_CARRYB_15__2_), .CI(u5_mult_82_SUMB_15__3_), .CO(
        u5_mult_82_CARRYB_16__2_), .S(u5_mult_82_SUMB_16__2_) );
  FA_X1 u5_mult_82_S2_16_1 ( .A(u5_mult_82_ab_16__1_), .B(
        u5_mult_82_CARRYB_15__1_), .CI(u5_mult_82_SUMB_15__2_), .CO(
        u5_mult_82_CARRYB_16__1_), .S(u5_mult_82_SUMB_16__1_) );
  FA_X1 u5_mult_82_S1_16_0 ( .A(u5_mult_82_ab_16__0_), .B(
        u5_mult_82_CARRYB_15__0_), .CI(u5_mult_82_SUMB_15__1_), .CO(
        u5_mult_82_CARRYB_16__0_), .S(u5_N16) );
  FA_X1 u5_mult_82_S3_17_51 ( .A(u5_mult_82_ab_17__51_), .B(
        u5_mult_82_CARRYB_16__51_), .CI(u5_mult_82_ab_16__52_), .CO(
        u5_mult_82_CARRYB_17__51_), .S(u5_mult_82_SUMB_17__51_) );
  FA_X1 u5_mult_82_S2_17_50 ( .A(u5_mult_82_ab_17__50_), .B(
        u5_mult_82_CARRYB_16__50_), .CI(u5_mult_82_SUMB_16__51_), .CO(
        u5_mult_82_CARRYB_17__50_), .S(u5_mult_82_SUMB_17__50_) );
  FA_X1 u5_mult_82_S2_17_49 ( .A(u5_mult_82_ab_17__49_), .B(
        u5_mult_82_CARRYB_16__49_), .CI(u5_mult_82_SUMB_16__50_), .CO(
        u5_mult_82_CARRYB_17__49_), .S(u5_mult_82_SUMB_17__49_) );
  FA_X1 u5_mult_82_S2_17_48 ( .A(u5_mult_82_ab_17__48_), .B(
        u5_mult_82_CARRYB_16__48_), .CI(u5_mult_82_SUMB_16__49_), .CO(
        u5_mult_82_CARRYB_17__48_), .S(u5_mult_82_SUMB_17__48_) );
  FA_X1 u5_mult_82_S2_17_47 ( .A(u5_mult_82_ab_17__47_), .B(
        u5_mult_82_CARRYB_16__47_), .CI(u5_mult_82_SUMB_16__48_), .CO(
        u5_mult_82_CARRYB_17__47_), .S(u5_mult_82_SUMB_17__47_) );
  FA_X1 u5_mult_82_S2_17_46 ( .A(u5_mult_82_ab_17__46_), .B(
        u5_mult_82_CARRYB_16__46_), .CI(u5_mult_82_SUMB_16__47_), .CO(
        u5_mult_82_CARRYB_17__46_), .S(u5_mult_82_SUMB_17__46_) );
  FA_X1 u5_mult_82_S2_17_45 ( .A(u5_mult_82_ab_17__45_), .B(
        u5_mult_82_CARRYB_16__45_), .CI(u5_mult_82_SUMB_16__46_), .CO(
        u5_mult_82_CARRYB_17__45_), .S(u5_mult_82_SUMB_17__45_) );
  FA_X1 u5_mult_82_S2_17_44 ( .A(u5_mult_82_ab_17__44_), .B(
        u5_mult_82_CARRYB_16__44_), .CI(u5_mult_82_SUMB_16__45_), .CO(
        u5_mult_82_CARRYB_17__44_), .S(u5_mult_82_SUMB_17__44_) );
  FA_X1 u5_mult_82_S2_17_43 ( .A(u5_mult_82_ab_17__43_), .B(
        u5_mult_82_CARRYB_16__43_), .CI(u5_mult_82_SUMB_16__44_), .CO(
        u5_mult_82_CARRYB_17__43_), .S(u5_mult_82_SUMB_17__43_) );
  FA_X1 u5_mult_82_S2_17_42 ( .A(u5_mult_82_ab_17__42_), .B(
        u5_mult_82_CARRYB_16__42_), .CI(u5_mult_82_SUMB_16__43_), .CO(
        u5_mult_82_CARRYB_17__42_), .S(u5_mult_82_SUMB_17__42_) );
  FA_X1 u5_mult_82_S2_17_41 ( .A(u5_mult_82_ab_17__41_), .B(
        u5_mult_82_CARRYB_16__41_), .CI(u5_mult_82_SUMB_16__42_), .CO(
        u5_mult_82_CARRYB_17__41_), .S(u5_mult_82_SUMB_17__41_) );
  FA_X1 u5_mult_82_S2_17_40 ( .A(u5_mult_82_ab_17__40_), .B(
        u5_mult_82_CARRYB_16__40_), .CI(u5_mult_82_SUMB_16__41_), .CO(
        u5_mult_82_CARRYB_17__40_), .S(u5_mult_82_SUMB_17__40_) );
  FA_X1 u5_mult_82_S2_17_39 ( .A(u5_mult_82_ab_17__39_), .B(
        u5_mult_82_CARRYB_16__39_), .CI(u5_mult_82_SUMB_16__40_), .CO(
        u5_mult_82_CARRYB_17__39_), .S(u5_mult_82_SUMB_17__39_) );
  FA_X1 u5_mult_82_S2_17_38 ( .A(u5_mult_82_ab_17__38_), .B(
        u5_mult_82_CARRYB_16__38_), .CI(u5_mult_82_SUMB_16__39_), .CO(
        u5_mult_82_CARRYB_17__38_), .S(u5_mult_82_SUMB_17__38_) );
  FA_X1 u5_mult_82_S2_17_37 ( .A(u5_mult_82_ab_17__37_), .B(
        u5_mult_82_CARRYB_16__37_), .CI(u5_mult_82_SUMB_16__38_), .CO(
        u5_mult_82_CARRYB_17__37_), .S(u5_mult_82_SUMB_17__37_) );
  FA_X1 u5_mult_82_S2_17_36 ( .A(u5_mult_82_ab_17__36_), .B(
        u5_mult_82_CARRYB_16__36_), .CI(u5_mult_82_SUMB_16__37_), .CO(
        u5_mult_82_CARRYB_17__36_), .S(u5_mult_82_SUMB_17__36_) );
  FA_X1 u5_mult_82_S2_17_35 ( .A(u5_mult_82_ab_17__35_), .B(
        u5_mult_82_CARRYB_16__35_), .CI(u5_mult_82_SUMB_16__36_), .CO(
        u5_mult_82_CARRYB_17__35_), .S(u5_mult_82_SUMB_17__35_) );
  FA_X1 u5_mult_82_S2_17_34 ( .A(u5_mult_82_ab_17__34_), .B(
        u5_mult_82_CARRYB_16__34_), .CI(u5_mult_82_SUMB_16__35_), .CO(
        u5_mult_82_CARRYB_17__34_), .S(u5_mult_82_SUMB_17__34_) );
  FA_X1 u5_mult_82_S2_17_33 ( .A(u5_mult_82_ab_17__33_), .B(
        u5_mult_82_CARRYB_16__33_), .CI(u5_mult_82_SUMB_16__34_), .CO(
        u5_mult_82_CARRYB_17__33_), .S(u5_mult_82_SUMB_17__33_) );
  FA_X1 u5_mult_82_S2_17_32 ( .A(u5_mult_82_ab_17__32_), .B(
        u5_mult_82_CARRYB_16__32_), .CI(u5_mult_82_SUMB_16__33_), .CO(
        u5_mult_82_CARRYB_17__32_), .S(u5_mult_82_SUMB_17__32_) );
  FA_X1 u5_mult_82_S2_17_31 ( .A(u5_mult_82_ab_17__31_), .B(
        u5_mult_82_CARRYB_16__31_), .CI(u5_mult_82_SUMB_16__32_), .CO(
        u5_mult_82_CARRYB_17__31_), .S(u5_mult_82_SUMB_17__31_) );
  FA_X1 u5_mult_82_S2_17_30 ( .A(u5_mult_82_ab_17__30_), .B(
        u5_mult_82_CARRYB_16__30_), .CI(u5_mult_82_SUMB_16__31_), .CO(
        u5_mult_82_CARRYB_17__30_), .S(u5_mult_82_SUMB_17__30_) );
  FA_X1 u5_mult_82_S2_17_29 ( .A(u5_mult_82_ab_17__29_), .B(
        u5_mult_82_CARRYB_16__29_), .CI(u5_mult_82_SUMB_16__30_), .CO(
        u5_mult_82_CARRYB_17__29_), .S(u5_mult_82_SUMB_17__29_) );
  FA_X1 u5_mult_82_S2_17_28 ( .A(u5_mult_82_ab_17__28_), .B(
        u5_mult_82_CARRYB_16__28_), .CI(u5_mult_82_SUMB_16__29_), .CO(
        u5_mult_82_CARRYB_17__28_), .S(u5_mult_82_SUMB_17__28_) );
  FA_X1 u5_mult_82_S2_17_27 ( .A(u5_mult_82_ab_17__27_), .B(
        u5_mult_82_CARRYB_16__27_), .CI(u5_mult_82_SUMB_16__28_), .CO(
        u5_mult_82_CARRYB_17__27_), .S(u5_mult_82_SUMB_17__27_) );
  FA_X1 u5_mult_82_S2_17_26 ( .A(u5_mult_82_ab_17__26_), .B(
        u5_mult_82_CARRYB_16__26_), .CI(u5_mult_82_SUMB_16__27_), .CO(
        u5_mult_82_CARRYB_17__26_), .S(u5_mult_82_SUMB_17__26_) );
  FA_X1 u5_mult_82_S2_17_25 ( .A(u5_mult_82_ab_17__25_), .B(
        u5_mult_82_CARRYB_16__25_), .CI(u5_mult_82_SUMB_16__26_), .CO(
        u5_mult_82_CARRYB_17__25_), .S(u5_mult_82_SUMB_17__25_) );
  FA_X1 u5_mult_82_S2_17_24 ( .A(u5_mult_82_ab_17__24_), .B(
        u5_mult_82_CARRYB_16__24_), .CI(u5_mult_82_SUMB_16__25_), .CO(
        u5_mult_82_CARRYB_17__24_), .S(u5_mult_82_SUMB_17__24_) );
  FA_X1 u5_mult_82_S2_17_23 ( .A(u5_mult_82_ab_17__23_), .B(
        u5_mult_82_CARRYB_16__23_), .CI(u5_mult_82_SUMB_16__24_), .CO(
        u5_mult_82_CARRYB_17__23_), .S(u5_mult_82_SUMB_17__23_) );
  FA_X1 u5_mult_82_S2_17_22 ( .A(u5_mult_82_ab_17__22_), .B(
        u5_mult_82_CARRYB_16__22_), .CI(u5_mult_82_SUMB_16__23_), .CO(
        u5_mult_82_CARRYB_17__22_), .S(u5_mult_82_SUMB_17__22_) );
  FA_X1 u5_mult_82_S2_17_21 ( .A(u5_mult_82_ab_17__21_), .B(
        u5_mult_82_CARRYB_16__21_), .CI(u5_mult_82_SUMB_16__22_), .CO(
        u5_mult_82_CARRYB_17__21_), .S(u5_mult_82_SUMB_17__21_) );
  FA_X1 u5_mult_82_S2_17_20 ( .A(u5_mult_82_ab_17__20_), .B(
        u5_mult_82_CARRYB_16__20_), .CI(u5_mult_82_SUMB_16__21_), .CO(
        u5_mult_82_CARRYB_17__20_), .S(u5_mult_82_SUMB_17__20_) );
  FA_X1 u5_mult_82_S2_17_19 ( .A(u5_mult_82_ab_17__19_), .B(
        u5_mult_82_CARRYB_16__19_), .CI(u5_mult_82_SUMB_16__20_), .CO(
        u5_mult_82_CARRYB_17__19_), .S(u5_mult_82_SUMB_17__19_) );
  FA_X1 u5_mult_82_S2_17_18 ( .A(u5_mult_82_ab_17__18_), .B(
        u5_mult_82_CARRYB_16__18_), .CI(u5_mult_82_SUMB_16__19_), .CO(
        u5_mult_82_CARRYB_17__18_), .S(u5_mult_82_SUMB_17__18_) );
  FA_X1 u5_mult_82_S2_17_17 ( .A(u5_mult_82_ab_17__17_), .B(
        u5_mult_82_CARRYB_16__17_), .CI(u5_mult_82_SUMB_16__18_), .CO(
        u5_mult_82_CARRYB_17__17_), .S(u5_mult_82_SUMB_17__17_) );
  FA_X1 u5_mult_82_S2_17_16 ( .A(u5_mult_82_ab_17__16_), .B(
        u5_mult_82_CARRYB_16__16_), .CI(u5_mult_82_SUMB_16__17_), .CO(
        u5_mult_82_CARRYB_17__16_), .S(u5_mult_82_SUMB_17__16_) );
  FA_X1 u5_mult_82_S2_17_15 ( .A(u5_mult_82_ab_17__15_), .B(
        u5_mult_82_CARRYB_16__15_), .CI(u5_mult_82_SUMB_16__16_), .CO(
        u5_mult_82_CARRYB_17__15_), .S(u5_mult_82_SUMB_17__15_) );
  FA_X1 u5_mult_82_S2_17_14 ( .A(u5_mult_82_ab_17__14_), .B(
        u5_mult_82_CARRYB_16__14_), .CI(u5_mult_82_SUMB_16__15_), .CO(
        u5_mult_82_CARRYB_17__14_), .S(u5_mult_82_SUMB_17__14_) );
  FA_X1 u5_mult_82_S2_17_13 ( .A(u5_mult_82_ab_17__13_), .B(
        u5_mult_82_CARRYB_16__13_), .CI(u5_mult_82_SUMB_16__14_), .CO(
        u5_mult_82_CARRYB_17__13_), .S(u5_mult_82_SUMB_17__13_) );
  FA_X1 u5_mult_82_S2_17_12 ( .A(u5_mult_82_ab_17__12_), .B(
        u5_mult_82_CARRYB_16__12_), .CI(u5_mult_82_SUMB_16__13_), .CO(
        u5_mult_82_CARRYB_17__12_), .S(u5_mult_82_SUMB_17__12_) );
  FA_X1 u5_mult_82_S2_17_11 ( .A(u5_mult_82_ab_17__11_), .B(
        u5_mult_82_CARRYB_16__11_), .CI(u5_mult_82_SUMB_16__12_), .CO(
        u5_mult_82_CARRYB_17__11_), .S(u5_mult_82_SUMB_17__11_) );
  FA_X1 u5_mult_82_S2_17_10 ( .A(u5_mult_82_ab_17__10_), .B(
        u5_mult_82_CARRYB_16__10_), .CI(u5_mult_82_SUMB_16__11_), .CO(
        u5_mult_82_CARRYB_17__10_), .S(u5_mult_82_SUMB_17__10_) );
  FA_X1 u5_mult_82_S2_17_9 ( .A(u5_mult_82_ab_17__9_), .B(
        u5_mult_82_CARRYB_16__9_), .CI(u5_mult_82_SUMB_16__10_), .CO(
        u5_mult_82_CARRYB_17__9_), .S(u5_mult_82_SUMB_17__9_) );
  FA_X1 u5_mult_82_S2_17_8 ( .A(u5_mult_82_ab_17__8_), .B(
        u5_mult_82_CARRYB_16__8_), .CI(u5_mult_82_SUMB_16__9_), .CO(
        u5_mult_82_CARRYB_17__8_), .S(u5_mult_82_SUMB_17__8_) );
  FA_X1 u5_mult_82_S2_17_7 ( .A(u5_mult_82_ab_17__7_), .B(
        u5_mult_82_CARRYB_16__7_), .CI(u5_mult_82_SUMB_16__8_), .CO(
        u5_mult_82_CARRYB_17__7_), .S(u5_mult_82_SUMB_17__7_) );
  FA_X1 u5_mult_82_S2_17_6 ( .A(u5_mult_82_ab_17__6_), .B(
        u5_mult_82_CARRYB_16__6_), .CI(u5_mult_82_SUMB_16__7_), .CO(
        u5_mult_82_CARRYB_17__6_), .S(u5_mult_82_SUMB_17__6_) );
  FA_X1 u5_mult_82_S2_17_5 ( .A(u5_mult_82_ab_17__5_), .B(
        u5_mult_82_CARRYB_16__5_), .CI(u5_mult_82_SUMB_16__6_), .CO(
        u5_mult_82_CARRYB_17__5_), .S(u5_mult_82_SUMB_17__5_) );
  FA_X1 u5_mult_82_S2_17_4 ( .A(u5_mult_82_ab_17__4_), .B(
        u5_mult_82_CARRYB_16__4_), .CI(u5_mult_82_SUMB_16__5_), .CO(
        u5_mult_82_CARRYB_17__4_), .S(u5_mult_82_SUMB_17__4_) );
  FA_X1 u5_mult_82_S2_17_3 ( .A(u5_mult_82_ab_17__3_), .B(
        u5_mult_82_CARRYB_16__3_), .CI(u5_mult_82_SUMB_16__4_), .CO(
        u5_mult_82_CARRYB_17__3_), .S(u5_mult_82_SUMB_17__3_) );
  FA_X1 u5_mult_82_S2_17_2 ( .A(u5_mult_82_ab_17__2_), .B(
        u5_mult_82_CARRYB_16__2_), .CI(u5_mult_82_SUMB_16__3_), .CO(
        u5_mult_82_CARRYB_17__2_), .S(u5_mult_82_SUMB_17__2_) );
  FA_X1 u5_mult_82_S2_17_1 ( .A(u5_mult_82_ab_17__1_), .B(
        u5_mult_82_CARRYB_16__1_), .CI(u5_mult_82_SUMB_16__2_), .CO(
        u5_mult_82_CARRYB_17__1_), .S(u5_mult_82_SUMB_17__1_) );
  FA_X1 u5_mult_82_S1_17_0 ( .A(u5_mult_82_ab_17__0_), .B(
        u5_mult_82_CARRYB_16__0_), .CI(u5_mult_82_SUMB_16__1_), .CO(
        u5_mult_82_CARRYB_17__0_), .S(u5_N17) );
  FA_X1 u5_mult_82_S3_18_51 ( .A(u5_mult_82_ab_18__51_), .B(
        u5_mult_82_CARRYB_17__51_), .CI(u5_mult_82_ab_17__52_), .CO(
        u5_mult_82_CARRYB_18__51_), .S(u5_mult_82_SUMB_18__51_) );
  FA_X1 u5_mult_82_S2_18_50 ( .A(u5_mult_82_ab_18__50_), .B(
        u5_mult_82_CARRYB_17__50_), .CI(u5_mult_82_SUMB_17__51_), .CO(
        u5_mult_82_CARRYB_18__50_), .S(u5_mult_82_SUMB_18__50_) );
  FA_X1 u5_mult_82_S2_18_49 ( .A(u5_mult_82_ab_18__49_), .B(
        u5_mult_82_CARRYB_17__49_), .CI(u5_mult_82_SUMB_17__50_), .CO(
        u5_mult_82_CARRYB_18__49_), .S(u5_mult_82_SUMB_18__49_) );
  FA_X1 u5_mult_82_S2_18_48 ( .A(u5_mult_82_ab_18__48_), .B(
        u5_mult_82_CARRYB_17__48_), .CI(u5_mult_82_SUMB_17__49_), .CO(
        u5_mult_82_CARRYB_18__48_), .S(u5_mult_82_SUMB_18__48_) );
  FA_X1 u5_mult_82_S2_18_47 ( .A(u5_mult_82_ab_18__47_), .B(
        u5_mult_82_CARRYB_17__47_), .CI(u5_mult_82_SUMB_17__48_), .CO(
        u5_mult_82_CARRYB_18__47_), .S(u5_mult_82_SUMB_18__47_) );
  FA_X1 u5_mult_82_S2_18_46 ( .A(u5_mult_82_ab_18__46_), .B(
        u5_mult_82_CARRYB_17__46_), .CI(u5_mult_82_SUMB_17__47_), .CO(
        u5_mult_82_CARRYB_18__46_), .S(u5_mult_82_SUMB_18__46_) );
  FA_X1 u5_mult_82_S2_18_45 ( .A(u5_mult_82_ab_18__45_), .B(
        u5_mult_82_CARRYB_17__45_), .CI(u5_mult_82_SUMB_17__46_), .CO(
        u5_mult_82_CARRYB_18__45_), .S(u5_mult_82_SUMB_18__45_) );
  FA_X1 u5_mult_82_S2_18_44 ( .A(u5_mult_82_ab_18__44_), .B(
        u5_mult_82_CARRYB_17__44_), .CI(u5_mult_82_SUMB_17__45_), .CO(
        u5_mult_82_CARRYB_18__44_), .S(u5_mult_82_SUMB_18__44_) );
  FA_X1 u5_mult_82_S2_18_43 ( .A(u5_mult_82_ab_18__43_), .B(
        u5_mult_82_CARRYB_17__43_), .CI(u5_mult_82_SUMB_17__44_), .CO(
        u5_mult_82_CARRYB_18__43_), .S(u5_mult_82_SUMB_18__43_) );
  FA_X1 u5_mult_82_S2_18_42 ( .A(u5_mult_82_ab_18__42_), .B(
        u5_mult_82_CARRYB_17__42_), .CI(u5_mult_82_SUMB_17__43_), .CO(
        u5_mult_82_CARRYB_18__42_), .S(u5_mult_82_SUMB_18__42_) );
  FA_X1 u5_mult_82_S2_18_41 ( .A(u5_mult_82_ab_18__41_), .B(
        u5_mult_82_CARRYB_17__41_), .CI(u5_mult_82_SUMB_17__42_), .CO(
        u5_mult_82_CARRYB_18__41_), .S(u5_mult_82_SUMB_18__41_) );
  FA_X1 u5_mult_82_S2_18_40 ( .A(u5_mult_82_ab_18__40_), .B(
        u5_mult_82_CARRYB_17__40_), .CI(u5_mult_82_SUMB_17__41_), .CO(
        u5_mult_82_CARRYB_18__40_), .S(u5_mult_82_SUMB_18__40_) );
  FA_X1 u5_mult_82_S2_18_39 ( .A(u5_mult_82_ab_18__39_), .B(
        u5_mult_82_CARRYB_17__39_), .CI(u5_mult_82_SUMB_17__40_), .CO(
        u5_mult_82_CARRYB_18__39_), .S(u5_mult_82_SUMB_18__39_) );
  FA_X1 u5_mult_82_S2_18_38 ( .A(u5_mult_82_ab_18__38_), .B(
        u5_mult_82_CARRYB_17__38_), .CI(u5_mult_82_SUMB_17__39_), .CO(
        u5_mult_82_CARRYB_18__38_), .S(u5_mult_82_SUMB_18__38_) );
  FA_X1 u5_mult_82_S2_18_37 ( .A(u5_mult_82_ab_18__37_), .B(
        u5_mult_82_CARRYB_17__37_), .CI(u5_mult_82_SUMB_17__38_), .CO(
        u5_mult_82_CARRYB_18__37_), .S(u5_mult_82_SUMB_18__37_) );
  FA_X1 u5_mult_82_S2_18_36 ( .A(u5_mult_82_ab_18__36_), .B(
        u5_mult_82_CARRYB_17__36_), .CI(u5_mult_82_SUMB_17__37_), .CO(
        u5_mult_82_CARRYB_18__36_), .S(u5_mult_82_SUMB_18__36_) );
  FA_X1 u5_mult_82_S2_18_35 ( .A(u5_mult_82_ab_18__35_), .B(
        u5_mult_82_CARRYB_17__35_), .CI(u5_mult_82_SUMB_17__36_), .CO(
        u5_mult_82_CARRYB_18__35_), .S(u5_mult_82_SUMB_18__35_) );
  FA_X1 u5_mult_82_S2_18_34 ( .A(u5_mult_82_ab_18__34_), .B(
        u5_mult_82_CARRYB_17__34_), .CI(u5_mult_82_SUMB_17__35_), .CO(
        u5_mult_82_CARRYB_18__34_), .S(u5_mult_82_SUMB_18__34_) );
  FA_X1 u5_mult_82_S2_18_33 ( .A(u5_mult_82_ab_18__33_), .B(
        u5_mult_82_CARRYB_17__33_), .CI(u5_mult_82_SUMB_17__34_), .CO(
        u5_mult_82_CARRYB_18__33_), .S(u5_mult_82_SUMB_18__33_) );
  FA_X1 u5_mult_82_S2_18_32 ( .A(u5_mult_82_ab_18__32_), .B(
        u5_mult_82_CARRYB_17__32_), .CI(u5_mult_82_SUMB_17__33_), .CO(
        u5_mult_82_CARRYB_18__32_), .S(u5_mult_82_SUMB_18__32_) );
  FA_X1 u5_mult_82_S2_18_31 ( .A(u5_mult_82_ab_18__31_), .B(
        u5_mult_82_CARRYB_17__31_), .CI(u5_mult_82_SUMB_17__32_), .CO(
        u5_mult_82_CARRYB_18__31_), .S(u5_mult_82_SUMB_18__31_) );
  FA_X1 u5_mult_82_S2_18_30 ( .A(u5_mult_82_ab_18__30_), .B(
        u5_mult_82_CARRYB_17__30_), .CI(u5_mult_82_SUMB_17__31_), .CO(
        u5_mult_82_CARRYB_18__30_), .S(u5_mult_82_SUMB_18__30_) );
  FA_X1 u5_mult_82_S2_18_29 ( .A(u5_mult_82_ab_18__29_), .B(
        u5_mult_82_CARRYB_17__29_), .CI(u5_mult_82_SUMB_17__30_), .CO(
        u5_mult_82_CARRYB_18__29_), .S(u5_mult_82_SUMB_18__29_) );
  FA_X1 u5_mult_82_S2_18_28 ( .A(u5_mult_82_ab_18__28_), .B(
        u5_mult_82_CARRYB_17__28_), .CI(u5_mult_82_SUMB_17__29_), .CO(
        u5_mult_82_CARRYB_18__28_), .S(u5_mult_82_SUMB_18__28_) );
  FA_X1 u5_mult_82_S2_18_27 ( .A(u5_mult_82_ab_18__27_), .B(
        u5_mult_82_CARRYB_17__27_), .CI(u5_mult_82_SUMB_17__28_), .CO(
        u5_mult_82_CARRYB_18__27_), .S(u5_mult_82_SUMB_18__27_) );
  FA_X1 u5_mult_82_S2_18_26 ( .A(u5_mult_82_ab_18__26_), .B(
        u5_mult_82_CARRYB_17__26_), .CI(u5_mult_82_SUMB_17__27_), .CO(
        u5_mult_82_CARRYB_18__26_), .S(u5_mult_82_SUMB_18__26_) );
  FA_X1 u5_mult_82_S2_18_25 ( .A(u5_mult_82_ab_18__25_), .B(
        u5_mult_82_CARRYB_17__25_), .CI(u5_mult_82_SUMB_17__26_), .CO(
        u5_mult_82_CARRYB_18__25_), .S(u5_mult_82_SUMB_18__25_) );
  FA_X1 u5_mult_82_S2_18_24 ( .A(u5_mult_82_ab_18__24_), .B(
        u5_mult_82_CARRYB_17__24_), .CI(u5_mult_82_SUMB_17__25_), .CO(
        u5_mult_82_CARRYB_18__24_), .S(u5_mult_82_SUMB_18__24_) );
  FA_X1 u5_mult_82_S2_18_23 ( .A(u5_mult_82_ab_18__23_), .B(
        u5_mult_82_CARRYB_17__23_), .CI(u5_mult_82_SUMB_17__24_), .CO(
        u5_mult_82_CARRYB_18__23_), .S(u5_mult_82_SUMB_18__23_) );
  FA_X1 u5_mult_82_S2_18_22 ( .A(u5_mult_82_ab_18__22_), .B(
        u5_mult_82_CARRYB_17__22_), .CI(u5_mult_82_SUMB_17__23_), .CO(
        u5_mult_82_CARRYB_18__22_), .S(u5_mult_82_SUMB_18__22_) );
  FA_X1 u5_mult_82_S2_18_21 ( .A(u5_mult_82_ab_18__21_), .B(
        u5_mult_82_CARRYB_17__21_), .CI(u5_mult_82_SUMB_17__22_), .CO(
        u5_mult_82_CARRYB_18__21_), .S(u5_mult_82_SUMB_18__21_) );
  FA_X1 u5_mult_82_S2_18_20 ( .A(u5_mult_82_ab_18__20_), .B(
        u5_mult_82_CARRYB_17__20_), .CI(u5_mult_82_SUMB_17__21_), .CO(
        u5_mult_82_CARRYB_18__20_), .S(u5_mult_82_SUMB_18__20_) );
  FA_X1 u5_mult_82_S2_18_19 ( .A(u5_mult_82_ab_18__19_), .B(
        u5_mult_82_CARRYB_17__19_), .CI(u5_mult_82_SUMB_17__20_), .CO(
        u5_mult_82_CARRYB_18__19_), .S(u5_mult_82_SUMB_18__19_) );
  FA_X1 u5_mult_82_S2_18_18 ( .A(u5_mult_82_ab_18__18_), .B(
        u5_mult_82_CARRYB_17__18_), .CI(u5_mult_82_SUMB_17__19_), .CO(
        u5_mult_82_CARRYB_18__18_), .S(u5_mult_82_SUMB_18__18_) );
  FA_X1 u5_mult_82_S2_18_17 ( .A(u5_mult_82_ab_18__17_), .B(
        u5_mult_82_CARRYB_17__17_), .CI(u5_mult_82_SUMB_17__18_), .CO(
        u5_mult_82_CARRYB_18__17_), .S(u5_mult_82_SUMB_18__17_) );
  FA_X1 u5_mult_82_S2_18_16 ( .A(u5_mult_82_ab_18__16_), .B(
        u5_mult_82_CARRYB_17__16_), .CI(u5_mult_82_SUMB_17__17_), .CO(
        u5_mult_82_CARRYB_18__16_), .S(u5_mult_82_SUMB_18__16_) );
  FA_X1 u5_mult_82_S2_18_15 ( .A(u5_mult_82_ab_18__15_), .B(
        u5_mult_82_CARRYB_17__15_), .CI(u5_mult_82_SUMB_17__16_), .CO(
        u5_mult_82_CARRYB_18__15_), .S(u5_mult_82_SUMB_18__15_) );
  FA_X1 u5_mult_82_S2_18_14 ( .A(u5_mult_82_ab_18__14_), .B(
        u5_mult_82_CARRYB_17__14_), .CI(u5_mult_82_SUMB_17__15_), .CO(
        u5_mult_82_CARRYB_18__14_), .S(u5_mult_82_SUMB_18__14_) );
  FA_X1 u5_mult_82_S2_18_13 ( .A(u5_mult_82_ab_18__13_), .B(
        u5_mult_82_CARRYB_17__13_), .CI(u5_mult_82_SUMB_17__14_), .CO(
        u5_mult_82_CARRYB_18__13_), .S(u5_mult_82_SUMB_18__13_) );
  FA_X1 u5_mult_82_S2_18_12 ( .A(u5_mult_82_ab_18__12_), .B(
        u5_mult_82_CARRYB_17__12_), .CI(u5_mult_82_SUMB_17__13_), .CO(
        u5_mult_82_CARRYB_18__12_), .S(u5_mult_82_SUMB_18__12_) );
  FA_X1 u5_mult_82_S2_18_11 ( .A(u5_mult_82_ab_18__11_), .B(
        u5_mult_82_CARRYB_17__11_), .CI(u5_mult_82_SUMB_17__12_), .CO(
        u5_mult_82_CARRYB_18__11_), .S(u5_mult_82_SUMB_18__11_) );
  FA_X1 u5_mult_82_S2_18_10 ( .A(u5_mult_82_ab_18__10_), .B(
        u5_mult_82_CARRYB_17__10_), .CI(u5_mult_82_SUMB_17__11_), .CO(
        u5_mult_82_CARRYB_18__10_), .S(u5_mult_82_SUMB_18__10_) );
  FA_X1 u5_mult_82_S2_18_9 ( .A(u5_mult_82_ab_18__9_), .B(
        u5_mult_82_CARRYB_17__9_), .CI(u5_mult_82_SUMB_17__10_), .CO(
        u5_mult_82_CARRYB_18__9_), .S(u5_mult_82_SUMB_18__9_) );
  FA_X1 u5_mult_82_S2_18_8 ( .A(u5_mult_82_ab_18__8_), .B(
        u5_mult_82_CARRYB_17__8_), .CI(u5_mult_82_SUMB_17__9_), .CO(
        u5_mult_82_CARRYB_18__8_), .S(u5_mult_82_SUMB_18__8_) );
  FA_X1 u5_mult_82_S2_18_7 ( .A(u5_mult_82_ab_18__7_), .B(
        u5_mult_82_CARRYB_17__7_), .CI(u5_mult_82_SUMB_17__8_), .CO(
        u5_mult_82_CARRYB_18__7_), .S(u5_mult_82_SUMB_18__7_) );
  FA_X1 u5_mult_82_S2_18_6 ( .A(u5_mult_82_ab_18__6_), .B(
        u5_mult_82_CARRYB_17__6_), .CI(u5_mult_82_SUMB_17__7_), .CO(
        u5_mult_82_CARRYB_18__6_), .S(u5_mult_82_SUMB_18__6_) );
  FA_X1 u5_mult_82_S2_18_5 ( .A(u5_mult_82_ab_18__5_), .B(
        u5_mult_82_CARRYB_17__5_), .CI(u5_mult_82_SUMB_17__6_), .CO(
        u5_mult_82_CARRYB_18__5_), .S(u5_mult_82_SUMB_18__5_) );
  FA_X1 u5_mult_82_S2_18_4 ( .A(u5_mult_82_ab_18__4_), .B(
        u5_mult_82_CARRYB_17__4_), .CI(u5_mult_82_SUMB_17__5_), .CO(
        u5_mult_82_CARRYB_18__4_), .S(u5_mult_82_SUMB_18__4_) );
  FA_X1 u5_mult_82_S2_18_3 ( .A(u5_mult_82_ab_18__3_), .B(
        u5_mult_82_CARRYB_17__3_), .CI(u5_mult_82_SUMB_17__4_), .CO(
        u5_mult_82_CARRYB_18__3_), .S(u5_mult_82_SUMB_18__3_) );
  FA_X1 u5_mult_82_S2_18_2 ( .A(u5_mult_82_ab_18__2_), .B(
        u5_mult_82_CARRYB_17__2_), .CI(u5_mult_82_SUMB_17__3_), .CO(
        u5_mult_82_CARRYB_18__2_), .S(u5_mult_82_SUMB_18__2_) );
  FA_X1 u5_mult_82_S2_18_1 ( .A(u5_mult_82_ab_18__1_), .B(
        u5_mult_82_CARRYB_17__1_), .CI(u5_mult_82_SUMB_17__2_), .CO(
        u5_mult_82_CARRYB_18__1_), .S(u5_mult_82_SUMB_18__1_) );
  FA_X1 u5_mult_82_S1_18_0 ( .A(u5_mult_82_ab_18__0_), .B(
        u5_mult_82_CARRYB_17__0_), .CI(u5_mult_82_SUMB_17__1_), .CO(
        u5_mult_82_CARRYB_18__0_), .S(u5_N18) );
  FA_X1 u5_mult_82_S3_19_51 ( .A(u5_mult_82_ab_19__51_), .B(
        u5_mult_82_CARRYB_18__51_), .CI(u5_mult_82_ab_18__52_), .CO(
        u5_mult_82_CARRYB_19__51_), .S(u5_mult_82_SUMB_19__51_) );
  FA_X1 u5_mult_82_S2_19_50 ( .A(u5_mult_82_ab_19__50_), .B(
        u5_mult_82_CARRYB_18__50_), .CI(u5_mult_82_SUMB_18__51_), .CO(
        u5_mult_82_CARRYB_19__50_), .S(u5_mult_82_SUMB_19__50_) );
  FA_X1 u5_mult_82_S2_19_49 ( .A(u5_mult_82_ab_19__49_), .B(
        u5_mult_82_CARRYB_18__49_), .CI(u5_mult_82_SUMB_18__50_), .CO(
        u5_mult_82_CARRYB_19__49_), .S(u5_mult_82_SUMB_19__49_) );
  FA_X1 u5_mult_82_S2_19_48 ( .A(u5_mult_82_ab_19__48_), .B(
        u5_mult_82_CARRYB_18__48_), .CI(u5_mult_82_SUMB_18__49_), .CO(
        u5_mult_82_CARRYB_19__48_), .S(u5_mult_82_SUMB_19__48_) );
  FA_X1 u5_mult_82_S2_19_47 ( .A(u5_mult_82_ab_19__47_), .B(
        u5_mult_82_CARRYB_18__47_), .CI(u5_mult_82_SUMB_18__48_), .CO(
        u5_mult_82_CARRYB_19__47_), .S(u5_mult_82_SUMB_19__47_) );
  FA_X1 u5_mult_82_S2_19_46 ( .A(u5_mult_82_ab_19__46_), .B(
        u5_mult_82_CARRYB_18__46_), .CI(u5_mult_82_SUMB_18__47_), .CO(
        u5_mult_82_CARRYB_19__46_), .S(u5_mult_82_SUMB_19__46_) );
  FA_X1 u5_mult_82_S2_19_45 ( .A(u5_mult_82_ab_19__45_), .B(
        u5_mult_82_CARRYB_18__45_), .CI(u5_mult_82_SUMB_18__46_), .CO(
        u5_mult_82_CARRYB_19__45_), .S(u5_mult_82_SUMB_19__45_) );
  FA_X1 u5_mult_82_S2_19_44 ( .A(u5_mult_82_ab_19__44_), .B(
        u5_mult_82_CARRYB_18__44_), .CI(u5_mult_82_SUMB_18__45_), .CO(
        u5_mult_82_CARRYB_19__44_), .S(u5_mult_82_SUMB_19__44_) );
  FA_X1 u5_mult_82_S2_19_43 ( .A(u5_mult_82_ab_19__43_), .B(
        u5_mult_82_CARRYB_18__43_), .CI(u5_mult_82_SUMB_18__44_), .CO(
        u5_mult_82_CARRYB_19__43_), .S(u5_mult_82_SUMB_19__43_) );
  FA_X1 u5_mult_82_S2_19_42 ( .A(u5_mult_82_ab_19__42_), .B(
        u5_mult_82_CARRYB_18__42_), .CI(u5_mult_82_SUMB_18__43_), .CO(
        u5_mult_82_CARRYB_19__42_), .S(u5_mult_82_SUMB_19__42_) );
  FA_X1 u5_mult_82_S2_19_41 ( .A(u5_mult_82_ab_19__41_), .B(
        u5_mult_82_CARRYB_18__41_), .CI(u5_mult_82_SUMB_18__42_), .CO(
        u5_mult_82_CARRYB_19__41_), .S(u5_mult_82_SUMB_19__41_) );
  FA_X1 u5_mult_82_S2_19_40 ( .A(u5_mult_82_ab_19__40_), .B(
        u5_mult_82_CARRYB_18__40_), .CI(u5_mult_82_SUMB_18__41_), .CO(
        u5_mult_82_CARRYB_19__40_), .S(u5_mult_82_SUMB_19__40_) );
  FA_X1 u5_mult_82_S2_19_39 ( .A(u5_mult_82_ab_19__39_), .B(
        u5_mult_82_CARRYB_18__39_), .CI(u5_mult_82_SUMB_18__40_), .CO(
        u5_mult_82_CARRYB_19__39_), .S(u5_mult_82_SUMB_19__39_) );
  FA_X1 u5_mult_82_S2_19_38 ( .A(u5_mult_82_ab_19__38_), .B(
        u5_mult_82_CARRYB_18__38_), .CI(u5_mult_82_SUMB_18__39_), .CO(
        u5_mult_82_CARRYB_19__38_), .S(u5_mult_82_SUMB_19__38_) );
  FA_X1 u5_mult_82_S2_19_37 ( .A(u5_mult_82_ab_19__37_), .B(
        u5_mult_82_CARRYB_18__37_), .CI(u5_mult_82_SUMB_18__38_), .CO(
        u5_mult_82_CARRYB_19__37_), .S(u5_mult_82_SUMB_19__37_) );
  FA_X1 u5_mult_82_S2_19_36 ( .A(u5_mult_82_ab_19__36_), .B(
        u5_mult_82_CARRYB_18__36_), .CI(u5_mult_82_SUMB_18__37_), .CO(
        u5_mult_82_CARRYB_19__36_), .S(u5_mult_82_SUMB_19__36_) );
  FA_X1 u5_mult_82_S2_19_35 ( .A(u5_mult_82_ab_19__35_), .B(
        u5_mult_82_CARRYB_18__35_), .CI(u5_mult_82_SUMB_18__36_), .CO(
        u5_mult_82_CARRYB_19__35_), .S(u5_mult_82_SUMB_19__35_) );
  FA_X1 u5_mult_82_S2_19_34 ( .A(u5_mult_82_ab_19__34_), .B(
        u5_mult_82_CARRYB_18__34_), .CI(u5_mult_82_SUMB_18__35_), .CO(
        u5_mult_82_CARRYB_19__34_), .S(u5_mult_82_SUMB_19__34_) );
  FA_X1 u5_mult_82_S2_19_33 ( .A(u5_mult_82_ab_19__33_), .B(
        u5_mult_82_CARRYB_18__33_), .CI(u5_mult_82_SUMB_18__34_), .CO(
        u5_mult_82_CARRYB_19__33_), .S(u5_mult_82_SUMB_19__33_) );
  FA_X1 u5_mult_82_S2_19_32 ( .A(u5_mult_82_ab_19__32_), .B(
        u5_mult_82_CARRYB_18__32_), .CI(u5_mult_82_SUMB_18__33_), .CO(
        u5_mult_82_CARRYB_19__32_), .S(u5_mult_82_SUMB_19__32_) );
  FA_X1 u5_mult_82_S2_19_31 ( .A(u5_mult_82_ab_19__31_), .B(
        u5_mult_82_CARRYB_18__31_), .CI(u5_mult_82_SUMB_18__32_), .CO(
        u5_mult_82_CARRYB_19__31_), .S(u5_mult_82_SUMB_19__31_) );
  FA_X1 u5_mult_82_S2_19_30 ( .A(u5_mult_82_ab_19__30_), .B(
        u5_mult_82_CARRYB_18__30_), .CI(u5_mult_82_SUMB_18__31_), .CO(
        u5_mult_82_CARRYB_19__30_), .S(u5_mult_82_SUMB_19__30_) );
  FA_X1 u5_mult_82_S2_19_29 ( .A(u5_mult_82_ab_19__29_), .B(
        u5_mult_82_CARRYB_18__29_), .CI(u5_mult_82_SUMB_18__30_), .CO(
        u5_mult_82_CARRYB_19__29_), .S(u5_mult_82_SUMB_19__29_) );
  FA_X1 u5_mult_82_S2_19_28 ( .A(u5_mult_82_ab_19__28_), .B(
        u5_mult_82_CARRYB_18__28_), .CI(u5_mult_82_SUMB_18__29_), .CO(
        u5_mult_82_CARRYB_19__28_), .S(u5_mult_82_SUMB_19__28_) );
  FA_X1 u5_mult_82_S2_19_27 ( .A(u5_mult_82_ab_19__27_), .B(
        u5_mult_82_CARRYB_18__27_), .CI(u5_mult_82_SUMB_18__28_), .CO(
        u5_mult_82_CARRYB_19__27_), .S(u5_mult_82_SUMB_19__27_) );
  FA_X1 u5_mult_82_S2_19_26 ( .A(u5_mult_82_ab_19__26_), .B(
        u5_mult_82_CARRYB_18__26_), .CI(u5_mult_82_SUMB_18__27_), .CO(
        u5_mult_82_CARRYB_19__26_), .S(u5_mult_82_SUMB_19__26_) );
  FA_X1 u5_mult_82_S2_19_25 ( .A(u5_mult_82_ab_19__25_), .B(
        u5_mult_82_CARRYB_18__25_), .CI(u5_mult_82_SUMB_18__26_), .CO(
        u5_mult_82_CARRYB_19__25_), .S(u5_mult_82_SUMB_19__25_) );
  FA_X1 u5_mult_82_S2_19_24 ( .A(u5_mult_82_ab_19__24_), .B(
        u5_mult_82_CARRYB_18__24_), .CI(u5_mult_82_SUMB_18__25_), .CO(
        u5_mult_82_CARRYB_19__24_), .S(u5_mult_82_SUMB_19__24_) );
  FA_X1 u5_mult_82_S2_19_23 ( .A(u5_mult_82_ab_19__23_), .B(
        u5_mult_82_CARRYB_18__23_), .CI(u5_mult_82_SUMB_18__24_), .CO(
        u5_mult_82_CARRYB_19__23_), .S(u5_mult_82_SUMB_19__23_) );
  FA_X1 u5_mult_82_S2_19_22 ( .A(u5_mult_82_ab_19__22_), .B(
        u5_mult_82_CARRYB_18__22_), .CI(u5_mult_82_SUMB_18__23_), .CO(
        u5_mult_82_CARRYB_19__22_), .S(u5_mult_82_SUMB_19__22_) );
  FA_X1 u5_mult_82_S2_19_21 ( .A(u5_mult_82_ab_19__21_), .B(
        u5_mult_82_CARRYB_18__21_), .CI(u5_mult_82_SUMB_18__22_), .CO(
        u5_mult_82_CARRYB_19__21_), .S(u5_mult_82_SUMB_19__21_) );
  FA_X1 u5_mult_82_S2_19_20 ( .A(u5_mult_82_ab_19__20_), .B(
        u5_mult_82_CARRYB_18__20_), .CI(u5_mult_82_SUMB_18__21_), .CO(
        u5_mult_82_CARRYB_19__20_), .S(u5_mult_82_SUMB_19__20_) );
  FA_X1 u5_mult_82_S2_19_19 ( .A(u5_mult_82_ab_19__19_), .B(
        u5_mult_82_CARRYB_18__19_), .CI(u5_mult_82_SUMB_18__20_), .CO(
        u5_mult_82_CARRYB_19__19_), .S(u5_mult_82_SUMB_19__19_) );
  FA_X1 u5_mult_82_S2_19_18 ( .A(u5_mult_82_ab_19__18_), .B(
        u5_mult_82_CARRYB_18__18_), .CI(u5_mult_82_SUMB_18__19_), .CO(
        u5_mult_82_CARRYB_19__18_), .S(u5_mult_82_SUMB_19__18_) );
  FA_X1 u5_mult_82_S2_19_17 ( .A(u5_mult_82_ab_19__17_), .B(
        u5_mult_82_CARRYB_18__17_), .CI(u5_mult_82_SUMB_18__18_), .CO(
        u5_mult_82_CARRYB_19__17_), .S(u5_mult_82_SUMB_19__17_) );
  FA_X1 u5_mult_82_S2_19_16 ( .A(u5_mult_82_ab_19__16_), .B(
        u5_mult_82_CARRYB_18__16_), .CI(u5_mult_82_SUMB_18__17_), .CO(
        u5_mult_82_CARRYB_19__16_), .S(u5_mult_82_SUMB_19__16_) );
  FA_X1 u5_mult_82_S2_19_15 ( .A(u5_mult_82_ab_19__15_), .B(
        u5_mult_82_CARRYB_18__15_), .CI(u5_mult_82_SUMB_18__16_), .CO(
        u5_mult_82_CARRYB_19__15_), .S(u5_mult_82_SUMB_19__15_) );
  FA_X1 u5_mult_82_S2_19_14 ( .A(u5_mult_82_ab_19__14_), .B(
        u5_mult_82_CARRYB_18__14_), .CI(u5_mult_82_SUMB_18__15_), .CO(
        u5_mult_82_CARRYB_19__14_), .S(u5_mult_82_SUMB_19__14_) );
  FA_X1 u5_mult_82_S2_19_13 ( .A(u5_mult_82_ab_19__13_), .B(
        u5_mult_82_CARRYB_18__13_), .CI(u5_mult_82_SUMB_18__14_), .CO(
        u5_mult_82_CARRYB_19__13_), .S(u5_mult_82_SUMB_19__13_) );
  FA_X1 u5_mult_82_S2_19_12 ( .A(u5_mult_82_ab_19__12_), .B(
        u5_mult_82_CARRYB_18__12_), .CI(u5_mult_82_SUMB_18__13_), .CO(
        u5_mult_82_CARRYB_19__12_), .S(u5_mult_82_SUMB_19__12_) );
  FA_X1 u5_mult_82_S2_19_11 ( .A(u5_mult_82_ab_19__11_), .B(
        u5_mult_82_CARRYB_18__11_), .CI(u5_mult_82_SUMB_18__12_), .CO(
        u5_mult_82_CARRYB_19__11_), .S(u5_mult_82_SUMB_19__11_) );
  FA_X1 u5_mult_82_S2_19_10 ( .A(u5_mult_82_ab_19__10_), .B(
        u5_mult_82_CARRYB_18__10_), .CI(u5_mult_82_SUMB_18__11_), .CO(
        u5_mult_82_CARRYB_19__10_), .S(u5_mult_82_SUMB_19__10_) );
  FA_X1 u5_mult_82_S2_19_9 ( .A(u5_mult_82_ab_19__9_), .B(
        u5_mult_82_CARRYB_18__9_), .CI(u5_mult_82_SUMB_18__10_), .CO(
        u5_mult_82_CARRYB_19__9_), .S(u5_mult_82_SUMB_19__9_) );
  FA_X1 u5_mult_82_S2_19_8 ( .A(u5_mult_82_ab_19__8_), .B(
        u5_mult_82_CARRYB_18__8_), .CI(u5_mult_82_SUMB_18__9_), .CO(
        u5_mult_82_CARRYB_19__8_), .S(u5_mult_82_SUMB_19__8_) );
  FA_X1 u5_mult_82_S2_19_7 ( .A(u5_mult_82_ab_19__7_), .B(
        u5_mult_82_CARRYB_18__7_), .CI(u5_mult_82_SUMB_18__8_), .CO(
        u5_mult_82_CARRYB_19__7_), .S(u5_mult_82_SUMB_19__7_) );
  FA_X1 u5_mult_82_S2_19_6 ( .A(u5_mult_82_ab_19__6_), .B(
        u5_mult_82_CARRYB_18__6_), .CI(u5_mult_82_SUMB_18__7_), .CO(
        u5_mult_82_CARRYB_19__6_), .S(u5_mult_82_SUMB_19__6_) );
  FA_X1 u5_mult_82_S2_19_5 ( .A(u5_mult_82_ab_19__5_), .B(
        u5_mult_82_CARRYB_18__5_), .CI(u5_mult_82_SUMB_18__6_), .CO(
        u5_mult_82_CARRYB_19__5_), .S(u5_mult_82_SUMB_19__5_) );
  FA_X1 u5_mult_82_S2_19_4 ( .A(u5_mult_82_ab_19__4_), .B(
        u5_mult_82_CARRYB_18__4_), .CI(u5_mult_82_SUMB_18__5_), .CO(
        u5_mult_82_CARRYB_19__4_), .S(u5_mult_82_SUMB_19__4_) );
  FA_X1 u5_mult_82_S2_19_3 ( .A(u5_mult_82_ab_19__3_), .B(
        u5_mult_82_CARRYB_18__3_), .CI(u5_mult_82_SUMB_18__4_), .CO(
        u5_mult_82_CARRYB_19__3_), .S(u5_mult_82_SUMB_19__3_) );
  FA_X1 u5_mult_82_S2_19_2 ( .A(u5_mult_82_ab_19__2_), .B(
        u5_mult_82_CARRYB_18__2_), .CI(u5_mult_82_SUMB_18__3_), .CO(
        u5_mult_82_CARRYB_19__2_), .S(u5_mult_82_SUMB_19__2_) );
  FA_X1 u5_mult_82_S2_19_1 ( .A(u5_mult_82_ab_19__1_), .B(
        u5_mult_82_CARRYB_18__1_), .CI(u5_mult_82_SUMB_18__2_), .CO(
        u5_mult_82_CARRYB_19__1_), .S(u5_mult_82_SUMB_19__1_) );
  FA_X1 u5_mult_82_S1_19_0 ( .A(u5_mult_82_ab_19__0_), .B(
        u5_mult_82_CARRYB_18__0_), .CI(u5_mult_82_SUMB_18__1_), .CO(
        u5_mult_82_CARRYB_19__0_), .S(u5_N19) );
  FA_X1 u5_mult_82_S3_20_51 ( .A(u5_mult_82_ab_20__51_), .B(
        u5_mult_82_CARRYB_19__51_), .CI(u5_mult_82_ab_19__52_), .CO(
        u5_mult_82_CARRYB_20__51_), .S(u5_mult_82_SUMB_20__51_) );
  FA_X1 u5_mult_82_S2_20_50 ( .A(u5_mult_82_ab_20__50_), .B(
        u5_mult_82_CARRYB_19__50_), .CI(u5_mult_82_SUMB_19__51_), .CO(
        u5_mult_82_CARRYB_20__50_), .S(u5_mult_82_SUMB_20__50_) );
  FA_X1 u5_mult_82_S2_20_49 ( .A(u5_mult_82_ab_20__49_), .B(
        u5_mult_82_CARRYB_19__49_), .CI(u5_mult_82_SUMB_19__50_), .CO(
        u5_mult_82_CARRYB_20__49_), .S(u5_mult_82_SUMB_20__49_) );
  FA_X1 u5_mult_82_S2_20_48 ( .A(u5_mult_82_ab_20__48_), .B(
        u5_mult_82_CARRYB_19__48_), .CI(u5_mult_82_SUMB_19__49_), .CO(
        u5_mult_82_CARRYB_20__48_), .S(u5_mult_82_SUMB_20__48_) );
  FA_X1 u5_mult_82_S2_20_47 ( .A(u5_mult_82_ab_20__47_), .B(
        u5_mult_82_CARRYB_19__47_), .CI(u5_mult_82_SUMB_19__48_), .CO(
        u5_mult_82_CARRYB_20__47_), .S(u5_mult_82_SUMB_20__47_) );
  FA_X1 u5_mult_82_S2_20_46 ( .A(u5_mult_82_ab_20__46_), .B(
        u5_mult_82_CARRYB_19__46_), .CI(u5_mult_82_SUMB_19__47_), .CO(
        u5_mult_82_CARRYB_20__46_), .S(u5_mult_82_SUMB_20__46_) );
  FA_X1 u5_mult_82_S2_20_45 ( .A(u5_mult_82_ab_20__45_), .B(
        u5_mult_82_CARRYB_19__45_), .CI(u5_mult_82_SUMB_19__46_), .CO(
        u5_mult_82_CARRYB_20__45_), .S(u5_mult_82_SUMB_20__45_) );
  FA_X1 u5_mult_82_S2_20_44 ( .A(u5_mult_82_ab_20__44_), .B(
        u5_mult_82_CARRYB_19__44_), .CI(u5_mult_82_SUMB_19__45_), .CO(
        u5_mult_82_CARRYB_20__44_), .S(u5_mult_82_SUMB_20__44_) );
  FA_X1 u5_mult_82_S2_20_43 ( .A(u5_mult_82_ab_20__43_), .B(
        u5_mult_82_CARRYB_19__43_), .CI(u5_mult_82_SUMB_19__44_), .CO(
        u5_mult_82_CARRYB_20__43_), .S(u5_mult_82_SUMB_20__43_) );
  FA_X1 u5_mult_82_S2_20_42 ( .A(u5_mult_82_ab_20__42_), .B(
        u5_mult_82_CARRYB_19__42_), .CI(u5_mult_82_SUMB_19__43_), .CO(
        u5_mult_82_CARRYB_20__42_), .S(u5_mult_82_SUMB_20__42_) );
  FA_X1 u5_mult_82_S2_20_41 ( .A(u5_mult_82_ab_20__41_), .B(
        u5_mult_82_CARRYB_19__41_), .CI(u5_mult_82_SUMB_19__42_), .CO(
        u5_mult_82_CARRYB_20__41_), .S(u5_mult_82_SUMB_20__41_) );
  FA_X1 u5_mult_82_S2_20_40 ( .A(u5_mult_82_ab_20__40_), .B(
        u5_mult_82_CARRYB_19__40_), .CI(u5_mult_82_SUMB_19__41_), .CO(
        u5_mult_82_CARRYB_20__40_), .S(u5_mult_82_SUMB_20__40_) );
  FA_X1 u5_mult_82_S2_20_39 ( .A(u5_mult_82_ab_20__39_), .B(
        u5_mult_82_CARRYB_19__39_), .CI(u5_mult_82_SUMB_19__40_), .CO(
        u5_mult_82_CARRYB_20__39_), .S(u5_mult_82_SUMB_20__39_) );
  FA_X1 u5_mult_82_S2_20_38 ( .A(u5_mult_82_ab_20__38_), .B(
        u5_mult_82_CARRYB_19__38_), .CI(u5_mult_82_SUMB_19__39_), .CO(
        u5_mult_82_CARRYB_20__38_), .S(u5_mult_82_SUMB_20__38_) );
  FA_X1 u5_mult_82_S2_20_37 ( .A(u5_mult_82_ab_20__37_), .B(
        u5_mult_82_CARRYB_19__37_), .CI(u5_mult_82_SUMB_19__38_), .CO(
        u5_mult_82_CARRYB_20__37_), .S(u5_mult_82_SUMB_20__37_) );
  FA_X1 u5_mult_82_S2_20_36 ( .A(u5_mult_82_ab_20__36_), .B(
        u5_mult_82_CARRYB_19__36_), .CI(u5_mult_82_SUMB_19__37_), .CO(
        u5_mult_82_CARRYB_20__36_), .S(u5_mult_82_SUMB_20__36_) );
  FA_X1 u5_mult_82_S2_20_35 ( .A(u5_mult_82_ab_20__35_), .B(
        u5_mult_82_CARRYB_19__35_), .CI(u5_mult_82_SUMB_19__36_), .CO(
        u5_mult_82_CARRYB_20__35_), .S(u5_mult_82_SUMB_20__35_) );
  FA_X1 u5_mult_82_S2_20_34 ( .A(u5_mult_82_ab_20__34_), .B(
        u5_mult_82_CARRYB_19__34_), .CI(u5_mult_82_SUMB_19__35_), .CO(
        u5_mult_82_CARRYB_20__34_), .S(u5_mult_82_SUMB_20__34_) );
  FA_X1 u5_mult_82_S2_20_33 ( .A(u5_mult_82_ab_20__33_), .B(
        u5_mult_82_CARRYB_19__33_), .CI(u5_mult_82_SUMB_19__34_), .CO(
        u5_mult_82_CARRYB_20__33_), .S(u5_mult_82_SUMB_20__33_) );
  FA_X1 u5_mult_82_S2_20_32 ( .A(u5_mult_82_ab_20__32_), .B(
        u5_mult_82_CARRYB_19__32_), .CI(u5_mult_82_SUMB_19__33_), .CO(
        u5_mult_82_CARRYB_20__32_), .S(u5_mult_82_SUMB_20__32_) );
  FA_X1 u5_mult_82_S2_20_31 ( .A(u5_mult_82_ab_20__31_), .B(
        u5_mult_82_CARRYB_19__31_), .CI(u5_mult_82_SUMB_19__32_), .CO(
        u5_mult_82_CARRYB_20__31_), .S(u5_mult_82_SUMB_20__31_) );
  FA_X1 u5_mult_82_S2_20_30 ( .A(u5_mult_82_ab_20__30_), .B(
        u5_mult_82_CARRYB_19__30_), .CI(u5_mult_82_SUMB_19__31_), .CO(
        u5_mult_82_CARRYB_20__30_), .S(u5_mult_82_SUMB_20__30_) );
  FA_X1 u5_mult_82_S2_20_29 ( .A(u5_mult_82_ab_20__29_), .B(
        u5_mult_82_CARRYB_19__29_), .CI(u5_mult_82_SUMB_19__30_), .CO(
        u5_mult_82_CARRYB_20__29_), .S(u5_mult_82_SUMB_20__29_) );
  FA_X1 u5_mult_82_S2_20_28 ( .A(u5_mult_82_ab_20__28_), .B(
        u5_mult_82_CARRYB_19__28_), .CI(u5_mult_82_SUMB_19__29_), .CO(
        u5_mult_82_CARRYB_20__28_), .S(u5_mult_82_SUMB_20__28_) );
  FA_X1 u5_mult_82_S2_20_27 ( .A(u5_mult_82_ab_20__27_), .B(
        u5_mult_82_CARRYB_19__27_), .CI(u5_mult_82_SUMB_19__28_), .CO(
        u5_mult_82_CARRYB_20__27_), .S(u5_mult_82_SUMB_20__27_) );
  FA_X1 u5_mult_82_S2_20_26 ( .A(u5_mult_82_ab_20__26_), .B(
        u5_mult_82_CARRYB_19__26_), .CI(u5_mult_82_SUMB_19__27_), .CO(
        u5_mult_82_CARRYB_20__26_), .S(u5_mult_82_SUMB_20__26_) );
  FA_X1 u5_mult_82_S2_20_25 ( .A(u5_mult_82_ab_20__25_), .B(
        u5_mult_82_CARRYB_19__25_), .CI(u5_mult_82_SUMB_19__26_), .CO(
        u5_mult_82_CARRYB_20__25_), .S(u5_mult_82_SUMB_20__25_) );
  FA_X1 u5_mult_82_S2_20_24 ( .A(u5_mult_82_ab_20__24_), .B(
        u5_mult_82_CARRYB_19__24_), .CI(u5_mult_82_SUMB_19__25_), .CO(
        u5_mult_82_CARRYB_20__24_), .S(u5_mult_82_SUMB_20__24_) );
  FA_X1 u5_mult_82_S2_20_23 ( .A(u5_mult_82_ab_20__23_), .B(
        u5_mult_82_CARRYB_19__23_), .CI(u5_mult_82_SUMB_19__24_), .CO(
        u5_mult_82_CARRYB_20__23_), .S(u5_mult_82_SUMB_20__23_) );
  FA_X1 u5_mult_82_S2_20_22 ( .A(u5_mult_82_ab_20__22_), .B(
        u5_mult_82_CARRYB_19__22_), .CI(u5_mult_82_SUMB_19__23_), .CO(
        u5_mult_82_CARRYB_20__22_), .S(u5_mult_82_SUMB_20__22_) );
  FA_X1 u5_mult_82_S2_20_21 ( .A(u5_mult_82_ab_20__21_), .B(
        u5_mult_82_CARRYB_19__21_), .CI(u5_mult_82_SUMB_19__22_), .CO(
        u5_mult_82_CARRYB_20__21_), .S(u5_mult_82_SUMB_20__21_) );
  FA_X1 u5_mult_82_S2_20_20 ( .A(u5_mult_82_ab_20__20_), .B(
        u5_mult_82_CARRYB_19__20_), .CI(u5_mult_82_SUMB_19__21_), .CO(
        u5_mult_82_CARRYB_20__20_), .S(u5_mult_82_SUMB_20__20_) );
  FA_X1 u5_mult_82_S2_20_19 ( .A(u5_mult_82_ab_20__19_), .B(
        u5_mult_82_CARRYB_19__19_), .CI(u5_mult_82_SUMB_19__20_), .CO(
        u5_mult_82_CARRYB_20__19_), .S(u5_mult_82_SUMB_20__19_) );
  FA_X1 u5_mult_82_S2_20_18 ( .A(u5_mult_82_ab_20__18_), .B(
        u5_mult_82_CARRYB_19__18_), .CI(u5_mult_82_SUMB_19__19_), .CO(
        u5_mult_82_CARRYB_20__18_), .S(u5_mult_82_SUMB_20__18_) );
  FA_X1 u5_mult_82_S2_20_17 ( .A(u5_mult_82_ab_20__17_), .B(
        u5_mult_82_CARRYB_19__17_), .CI(u5_mult_82_SUMB_19__18_), .CO(
        u5_mult_82_CARRYB_20__17_), .S(u5_mult_82_SUMB_20__17_) );
  FA_X1 u5_mult_82_S2_20_16 ( .A(u5_mult_82_ab_20__16_), .B(
        u5_mult_82_CARRYB_19__16_), .CI(u5_mult_82_SUMB_19__17_), .CO(
        u5_mult_82_CARRYB_20__16_), .S(u5_mult_82_SUMB_20__16_) );
  FA_X1 u5_mult_82_S2_20_15 ( .A(u5_mult_82_ab_20__15_), .B(
        u5_mult_82_CARRYB_19__15_), .CI(u5_mult_82_SUMB_19__16_), .CO(
        u5_mult_82_CARRYB_20__15_), .S(u5_mult_82_SUMB_20__15_) );
  FA_X1 u5_mult_82_S2_20_14 ( .A(u5_mult_82_ab_20__14_), .B(
        u5_mult_82_CARRYB_19__14_), .CI(u5_mult_82_SUMB_19__15_), .CO(
        u5_mult_82_CARRYB_20__14_), .S(u5_mult_82_SUMB_20__14_) );
  FA_X1 u5_mult_82_S2_20_13 ( .A(u5_mult_82_ab_20__13_), .B(
        u5_mult_82_CARRYB_19__13_), .CI(u5_mult_82_SUMB_19__14_), .CO(
        u5_mult_82_CARRYB_20__13_), .S(u5_mult_82_SUMB_20__13_) );
  FA_X1 u5_mult_82_S2_20_12 ( .A(u5_mult_82_ab_20__12_), .B(
        u5_mult_82_CARRYB_19__12_), .CI(u5_mult_82_SUMB_19__13_), .CO(
        u5_mult_82_CARRYB_20__12_), .S(u5_mult_82_SUMB_20__12_) );
  FA_X1 u5_mult_82_S2_20_11 ( .A(u5_mult_82_ab_20__11_), .B(
        u5_mult_82_CARRYB_19__11_), .CI(u5_mult_82_SUMB_19__12_), .CO(
        u5_mult_82_CARRYB_20__11_), .S(u5_mult_82_SUMB_20__11_) );
  FA_X1 u5_mult_82_S2_20_10 ( .A(u5_mult_82_ab_20__10_), .B(
        u5_mult_82_CARRYB_19__10_), .CI(u5_mult_82_SUMB_19__11_), .CO(
        u5_mult_82_CARRYB_20__10_), .S(u5_mult_82_SUMB_20__10_) );
  FA_X1 u5_mult_82_S2_20_9 ( .A(u5_mult_82_ab_20__9_), .B(
        u5_mult_82_CARRYB_19__9_), .CI(u5_mult_82_SUMB_19__10_), .CO(
        u5_mult_82_CARRYB_20__9_), .S(u5_mult_82_SUMB_20__9_) );
  FA_X1 u5_mult_82_S2_20_8 ( .A(u5_mult_82_ab_20__8_), .B(
        u5_mult_82_CARRYB_19__8_), .CI(u5_mult_82_SUMB_19__9_), .CO(
        u5_mult_82_CARRYB_20__8_), .S(u5_mult_82_SUMB_20__8_) );
  FA_X1 u5_mult_82_S2_20_7 ( .A(u5_mult_82_ab_20__7_), .B(
        u5_mult_82_CARRYB_19__7_), .CI(u5_mult_82_SUMB_19__8_), .CO(
        u5_mult_82_CARRYB_20__7_), .S(u5_mult_82_SUMB_20__7_) );
  FA_X1 u5_mult_82_S2_20_6 ( .A(u5_mult_82_ab_20__6_), .B(
        u5_mult_82_CARRYB_19__6_), .CI(u5_mult_82_SUMB_19__7_), .CO(
        u5_mult_82_CARRYB_20__6_), .S(u5_mult_82_SUMB_20__6_) );
  FA_X1 u5_mult_82_S2_20_5 ( .A(u5_mult_82_ab_20__5_), .B(
        u5_mult_82_CARRYB_19__5_), .CI(u5_mult_82_SUMB_19__6_), .CO(
        u5_mult_82_CARRYB_20__5_), .S(u5_mult_82_SUMB_20__5_) );
  FA_X1 u5_mult_82_S2_20_4 ( .A(u5_mult_82_ab_20__4_), .B(
        u5_mult_82_CARRYB_19__4_), .CI(u5_mult_82_SUMB_19__5_), .CO(
        u5_mult_82_CARRYB_20__4_), .S(u5_mult_82_SUMB_20__4_) );
  FA_X1 u5_mult_82_S2_20_3 ( .A(u5_mult_82_ab_20__3_), .B(
        u5_mult_82_CARRYB_19__3_), .CI(u5_mult_82_SUMB_19__4_), .CO(
        u5_mult_82_CARRYB_20__3_), .S(u5_mult_82_SUMB_20__3_) );
  FA_X1 u5_mult_82_S2_20_2 ( .A(u5_mult_82_ab_20__2_), .B(
        u5_mult_82_CARRYB_19__2_), .CI(u5_mult_82_SUMB_19__3_), .CO(
        u5_mult_82_CARRYB_20__2_), .S(u5_mult_82_SUMB_20__2_) );
  FA_X1 u5_mult_82_S2_20_1 ( .A(u5_mult_82_ab_20__1_), .B(
        u5_mult_82_CARRYB_19__1_), .CI(u5_mult_82_SUMB_19__2_), .CO(
        u5_mult_82_CARRYB_20__1_), .S(u5_mult_82_SUMB_20__1_) );
  FA_X1 u5_mult_82_S1_20_0 ( .A(u5_mult_82_ab_20__0_), .B(
        u5_mult_82_CARRYB_19__0_), .CI(u5_mult_82_SUMB_19__1_), .CO(
        u5_mult_82_CARRYB_20__0_), .S(u5_N20) );
  FA_X1 u5_mult_82_S3_21_51 ( .A(u5_mult_82_ab_21__51_), .B(
        u5_mult_82_CARRYB_20__51_), .CI(u5_mult_82_ab_20__52_), .CO(
        u5_mult_82_CARRYB_21__51_), .S(u5_mult_82_SUMB_21__51_) );
  FA_X1 u5_mult_82_S2_21_50 ( .A(u5_mult_82_ab_21__50_), .B(
        u5_mult_82_CARRYB_20__50_), .CI(u5_mult_82_SUMB_20__51_), .CO(
        u5_mult_82_CARRYB_21__50_), .S(u5_mult_82_SUMB_21__50_) );
  FA_X1 u5_mult_82_S2_21_49 ( .A(u5_mult_82_ab_21__49_), .B(
        u5_mult_82_CARRYB_20__49_), .CI(u5_mult_82_SUMB_20__50_), .CO(
        u5_mult_82_CARRYB_21__49_), .S(u5_mult_82_SUMB_21__49_) );
  FA_X1 u5_mult_82_S2_21_48 ( .A(u5_mult_82_ab_21__48_), .B(
        u5_mult_82_CARRYB_20__48_), .CI(u5_mult_82_SUMB_20__49_), .CO(
        u5_mult_82_CARRYB_21__48_), .S(u5_mult_82_SUMB_21__48_) );
  FA_X1 u5_mult_82_S2_21_47 ( .A(u5_mult_82_ab_21__47_), .B(
        u5_mult_82_CARRYB_20__47_), .CI(u5_mult_82_SUMB_20__48_), .CO(
        u5_mult_82_CARRYB_21__47_), .S(u5_mult_82_SUMB_21__47_) );
  FA_X1 u5_mult_82_S2_21_46 ( .A(u5_mult_82_ab_21__46_), .B(
        u5_mult_82_CARRYB_20__46_), .CI(u5_mult_82_SUMB_20__47_), .CO(
        u5_mult_82_CARRYB_21__46_), .S(u5_mult_82_SUMB_21__46_) );
  FA_X1 u5_mult_82_S2_21_45 ( .A(u5_mult_82_ab_21__45_), .B(
        u5_mult_82_CARRYB_20__45_), .CI(u5_mult_82_SUMB_20__46_), .CO(
        u5_mult_82_CARRYB_21__45_), .S(u5_mult_82_SUMB_21__45_) );
  FA_X1 u5_mult_82_S2_21_44 ( .A(u5_mult_82_ab_21__44_), .B(
        u5_mult_82_CARRYB_20__44_), .CI(u5_mult_82_SUMB_20__45_), .CO(
        u5_mult_82_CARRYB_21__44_), .S(u5_mult_82_SUMB_21__44_) );
  FA_X1 u5_mult_82_S2_21_43 ( .A(u5_mult_82_ab_21__43_), .B(
        u5_mult_82_CARRYB_20__43_), .CI(u5_mult_82_SUMB_20__44_), .CO(
        u5_mult_82_CARRYB_21__43_), .S(u5_mult_82_SUMB_21__43_) );
  FA_X1 u5_mult_82_S2_21_42 ( .A(u5_mult_82_ab_21__42_), .B(
        u5_mult_82_CARRYB_20__42_), .CI(u5_mult_82_SUMB_20__43_), .CO(
        u5_mult_82_CARRYB_21__42_), .S(u5_mult_82_SUMB_21__42_) );
  FA_X1 u5_mult_82_S2_21_41 ( .A(u5_mult_82_ab_21__41_), .B(
        u5_mult_82_CARRYB_20__41_), .CI(u5_mult_82_SUMB_20__42_), .CO(
        u5_mult_82_CARRYB_21__41_), .S(u5_mult_82_SUMB_21__41_) );
  FA_X1 u5_mult_82_S2_21_40 ( .A(u5_mult_82_ab_21__40_), .B(
        u5_mult_82_CARRYB_20__40_), .CI(u5_mult_82_SUMB_20__41_), .CO(
        u5_mult_82_CARRYB_21__40_), .S(u5_mult_82_SUMB_21__40_) );
  FA_X1 u5_mult_82_S2_21_39 ( .A(u5_mult_82_ab_21__39_), .B(
        u5_mult_82_CARRYB_20__39_), .CI(u5_mult_82_SUMB_20__40_), .CO(
        u5_mult_82_CARRYB_21__39_), .S(u5_mult_82_SUMB_21__39_) );
  FA_X1 u5_mult_82_S2_21_38 ( .A(u5_mult_82_ab_21__38_), .B(
        u5_mult_82_CARRYB_20__38_), .CI(u5_mult_82_SUMB_20__39_), .CO(
        u5_mult_82_CARRYB_21__38_), .S(u5_mult_82_SUMB_21__38_) );
  FA_X1 u5_mult_82_S2_21_37 ( .A(u5_mult_82_ab_21__37_), .B(
        u5_mult_82_CARRYB_20__37_), .CI(u5_mult_82_SUMB_20__38_), .CO(
        u5_mult_82_CARRYB_21__37_), .S(u5_mult_82_SUMB_21__37_) );
  FA_X1 u5_mult_82_S2_21_36 ( .A(u5_mult_82_ab_21__36_), .B(
        u5_mult_82_CARRYB_20__36_), .CI(u5_mult_82_SUMB_20__37_), .CO(
        u5_mult_82_CARRYB_21__36_), .S(u5_mult_82_SUMB_21__36_) );
  FA_X1 u5_mult_82_S2_21_35 ( .A(u5_mult_82_ab_21__35_), .B(
        u5_mult_82_CARRYB_20__35_), .CI(u5_mult_82_SUMB_20__36_), .CO(
        u5_mult_82_CARRYB_21__35_), .S(u5_mult_82_SUMB_21__35_) );
  FA_X1 u5_mult_82_S2_21_34 ( .A(u5_mult_82_ab_21__34_), .B(
        u5_mult_82_CARRYB_20__34_), .CI(u5_mult_82_SUMB_20__35_), .CO(
        u5_mult_82_CARRYB_21__34_), .S(u5_mult_82_SUMB_21__34_) );
  FA_X1 u5_mult_82_S2_21_33 ( .A(u5_mult_82_ab_21__33_), .B(
        u5_mult_82_CARRYB_20__33_), .CI(u5_mult_82_SUMB_20__34_), .CO(
        u5_mult_82_CARRYB_21__33_), .S(u5_mult_82_SUMB_21__33_) );
  FA_X1 u5_mult_82_S2_21_32 ( .A(u5_mult_82_ab_21__32_), .B(
        u5_mult_82_CARRYB_20__32_), .CI(u5_mult_82_SUMB_20__33_), .CO(
        u5_mult_82_CARRYB_21__32_), .S(u5_mult_82_SUMB_21__32_) );
  FA_X1 u5_mult_82_S2_21_31 ( .A(u5_mult_82_ab_21__31_), .B(
        u5_mult_82_CARRYB_20__31_), .CI(u5_mult_82_SUMB_20__32_), .CO(
        u5_mult_82_CARRYB_21__31_), .S(u5_mult_82_SUMB_21__31_) );
  FA_X1 u5_mult_82_S2_21_30 ( .A(u5_mult_82_ab_21__30_), .B(
        u5_mult_82_CARRYB_20__30_), .CI(u5_mult_82_SUMB_20__31_), .CO(
        u5_mult_82_CARRYB_21__30_), .S(u5_mult_82_SUMB_21__30_) );
  FA_X1 u5_mult_82_S2_21_29 ( .A(u5_mult_82_ab_21__29_), .B(
        u5_mult_82_CARRYB_20__29_), .CI(u5_mult_82_SUMB_20__30_), .CO(
        u5_mult_82_CARRYB_21__29_), .S(u5_mult_82_SUMB_21__29_) );
  FA_X1 u5_mult_82_S2_21_28 ( .A(u5_mult_82_ab_21__28_), .B(
        u5_mult_82_CARRYB_20__28_), .CI(u5_mult_82_SUMB_20__29_), .CO(
        u5_mult_82_CARRYB_21__28_), .S(u5_mult_82_SUMB_21__28_) );
  FA_X1 u5_mult_82_S2_21_27 ( .A(u5_mult_82_ab_21__27_), .B(
        u5_mult_82_CARRYB_20__27_), .CI(u5_mult_82_SUMB_20__28_), .CO(
        u5_mult_82_CARRYB_21__27_), .S(u5_mult_82_SUMB_21__27_) );
  FA_X1 u5_mult_82_S2_21_26 ( .A(u5_mult_82_ab_21__26_), .B(
        u5_mult_82_CARRYB_20__26_), .CI(u5_mult_82_SUMB_20__27_), .CO(
        u5_mult_82_CARRYB_21__26_), .S(u5_mult_82_SUMB_21__26_) );
  FA_X1 u5_mult_82_S2_21_25 ( .A(u5_mult_82_ab_21__25_), .B(
        u5_mult_82_CARRYB_20__25_), .CI(u5_mult_82_SUMB_20__26_), .CO(
        u5_mult_82_CARRYB_21__25_), .S(u5_mult_82_SUMB_21__25_) );
  FA_X1 u5_mult_82_S2_21_24 ( .A(u5_mult_82_ab_21__24_), .B(
        u5_mult_82_CARRYB_20__24_), .CI(u5_mult_82_SUMB_20__25_), .CO(
        u5_mult_82_CARRYB_21__24_), .S(u5_mult_82_SUMB_21__24_) );
  FA_X1 u5_mult_82_S2_21_23 ( .A(u5_mult_82_ab_21__23_), .B(
        u5_mult_82_CARRYB_20__23_), .CI(u5_mult_82_SUMB_20__24_), .CO(
        u5_mult_82_CARRYB_21__23_), .S(u5_mult_82_SUMB_21__23_) );
  FA_X1 u5_mult_82_S2_21_22 ( .A(u5_mult_82_ab_21__22_), .B(
        u5_mult_82_CARRYB_20__22_), .CI(u5_mult_82_SUMB_20__23_), .CO(
        u5_mult_82_CARRYB_21__22_), .S(u5_mult_82_SUMB_21__22_) );
  FA_X1 u5_mult_82_S2_21_21 ( .A(u5_mult_82_ab_21__21_), .B(
        u5_mult_82_CARRYB_20__21_), .CI(u5_mult_82_SUMB_20__22_), .CO(
        u5_mult_82_CARRYB_21__21_), .S(u5_mult_82_SUMB_21__21_) );
  FA_X1 u5_mult_82_S2_21_20 ( .A(u5_mult_82_ab_21__20_), .B(
        u5_mult_82_CARRYB_20__20_), .CI(u5_mult_82_SUMB_20__21_), .CO(
        u5_mult_82_CARRYB_21__20_), .S(u5_mult_82_SUMB_21__20_) );
  FA_X1 u5_mult_82_S2_21_19 ( .A(u5_mult_82_ab_21__19_), .B(
        u5_mult_82_CARRYB_20__19_), .CI(u5_mult_82_SUMB_20__20_), .CO(
        u5_mult_82_CARRYB_21__19_), .S(u5_mult_82_SUMB_21__19_) );
  FA_X1 u5_mult_82_S2_21_18 ( .A(u5_mult_82_ab_21__18_), .B(
        u5_mult_82_CARRYB_20__18_), .CI(u5_mult_82_SUMB_20__19_), .CO(
        u5_mult_82_CARRYB_21__18_), .S(u5_mult_82_SUMB_21__18_) );
  FA_X1 u5_mult_82_S2_21_17 ( .A(u5_mult_82_ab_21__17_), .B(
        u5_mult_82_CARRYB_20__17_), .CI(u5_mult_82_SUMB_20__18_), .CO(
        u5_mult_82_CARRYB_21__17_), .S(u5_mult_82_SUMB_21__17_) );
  FA_X1 u5_mult_82_S2_21_16 ( .A(u5_mult_82_ab_21__16_), .B(
        u5_mult_82_CARRYB_20__16_), .CI(u5_mult_82_SUMB_20__17_), .CO(
        u5_mult_82_CARRYB_21__16_), .S(u5_mult_82_SUMB_21__16_) );
  FA_X1 u5_mult_82_S2_21_15 ( .A(u5_mult_82_ab_21__15_), .B(
        u5_mult_82_CARRYB_20__15_), .CI(u5_mult_82_SUMB_20__16_), .CO(
        u5_mult_82_CARRYB_21__15_), .S(u5_mult_82_SUMB_21__15_) );
  FA_X1 u5_mult_82_S2_21_14 ( .A(u5_mult_82_ab_21__14_), .B(
        u5_mult_82_CARRYB_20__14_), .CI(u5_mult_82_SUMB_20__15_), .CO(
        u5_mult_82_CARRYB_21__14_), .S(u5_mult_82_SUMB_21__14_) );
  FA_X1 u5_mult_82_S2_21_13 ( .A(u5_mult_82_ab_21__13_), .B(
        u5_mult_82_CARRYB_20__13_), .CI(u5_mult_82_SUMB_20__14_), .CO(
        u5_mult_82_CARRYB_21__13_), .S(u5_mult_82_SUMB_21__13_) );
  FA_X1 u5_mult_82_S2_21_12 ( .A(u5_mult_82_ab_21__12_), .B(
        u5_mult_82_CARRYB_20__12_), .CI(u5_mult_82_SUMB_20__13_), .CO(
        u5_mult_82_CARRYB_21__12_), .S(u5_mult_82_SUMB_21__12_) );
  FA_X1 u5_mult_82_S2_21_11 ( .A(u5_mult_82_ab_21__11_), .B(
        u5_mult_82_CARRYB_20__11_), .CI(u5_mult_82_SUMB_20__12_), .CO(
        u5_mult_82_CARRYB_21__11_), .S(u5_mult_82_SUMB_21__11_) );
  FA_X1 u5_mult_82_S2_21_10 ( .A(u5_mult_82_ab_21__10_), .B(
        u5_mult_82_CARRYB_20__10_), .CI(u5_mult_82_SUMB_20__11_), .CO(
        u5_mult_82_CARRYB_21__10_), .S(u5_mult_82_SUMB_21__10_) );
  FA_X1 u5_mult_82_S2_21_9 ( .A(u5_mult_82_ab_21__9_), .B(
        u5_mult_82_CARRYB_20__9_), .CI(u5_mult_82_SUMB_20__10_), .CO(
        u5_mult_82_CARRYB_21__9_), .S(u5_mult_82_SUMB_21__9_) );
  FA_X1 u5_mult_82_S2_21_8 ( .A(u5_mult_82_ab_21__8_), .B(
        u5_mult_82_CARRYB_20__8_), .CI(u5_mult_82_SUMB_20__9_), .CO(
        u5_mult_82_CARRYB_21__8_), .S(u5_mult_82_SUMB_21__8_) );
  FA_X1 u5_mult_82_S2_21_7 ( .A(u5_mult_82_ab_21__7_), .B(
        u5_mult_82_CARRYB_20__7_), .CI(u5_mult_82_SUMB_20__8_), .CO(
        u5_mult_82_CARRYB_21__7_), .S(u5_mult_82_SUMB_21__7_) );
  FA_X1 u5_mult_82_S2_21_6 ( .A(u5_mult_82_ab_21__6_), .B(
        u5_mult_82_CARRYB_20__6_), .CI(u5_mult_82_SUMB_20__7_), .CO(
        u5_mult_82_CARRYB_21__6_), .S(u5_mult_82_SUMB_21__6_) );
  FA_X1 u5_mult_82_S2_21_5 ( .A(u5_mult_82_ab_21__5_), .B(
        u5_mult_82_CARRYB_20__5_), .CI(u5_mult_82_SUMB_20__6_), .CO(
        u5_mult_82_CARRYB_21__5_), .S(u5_mult_82_SUMB_21__5_) );
  FA_X1 u5_mult_82_S2_21_4 ( .A(u5_mult_82_ab_21__4_), .B(
        u5_mult_82_CARRYB_20__4_), .CI(u5_mult_82_SUMB_20__5_), .CO(
        u5_mult_82_CARRYB_21__4_), .S(u5_mult_82_SUMB_21__4_) );
  FA_X1 u5_mult_82_S2_21_3 ( .A(u5_mult_82_ab_21__3_), .B(
        u5_mult_82_CARRYB_20__3_), .CI(u5_mult_82_SUMB_20__4_), .CO(
        u5_mult_82_CARRYB_21__3_), .S(u5_mult_82_SUMB_21__3_) );
  FA_X1 u5_mult_82_S2_21_2 ( .A(u5_mult_82_ab_21__2_), .B(
        u5_mult_82_CARRYB_20__2_), .CI(u5_mult_82_SUMB_20__3_), .CO(
        u5_mult_82_CARRYB_21__2_), .S(u5_mult_82_SUMB_21__2_) );
  FA_X1 u5_mult_82_S2_21_1 ( .A(u5_mult_82_ab_21__1_), .B(
        u5_mult_82_CARRYB_20__1_), .CI(u5_mult_82_SUMB_20__2_), .CO(
        u5_mult_82_CARRYB_21__1_), .S(u5_mult_82_SUMB_21__1_) );
  FA_X1 u5_mult_82_S1_21_0 ( .A(u5_mult_82_ab_21__0_), .B(
        u5_mult_82_CARRYB_20__0_), .CI(u5_mult_82_SUMB_20__1_), .CO(
        u5_mult_82_CARRYB_21__0_), .S(u5_N21) );
  FA_X1 u5_mult_82_S3_22_51 ( .A(u5_mult_82_ab_22__51_), .B(
        u5_mult_82_CARRYB_21__51_), .CI(u5_mult_82_ab_21__52_), .CO(
        u5_mult_82_CARRYB_22__51_), .S(u5_mult_82_SUMB_22__51_) );
  FA_X1 u5_mult_82_S2_22_50 ( .A(u5_mult_82_ab_22__50_), .B(
        u5_mult_82_CARRYB_21__50_), .CI(u5_mult_82_SUMB_21__51_), .CO(
        u5_mult_82_CARRYB_22__50_), .S(u5_mult_82_SUMB_22__50_) );
  FA_X1 u5_mult_82_S2_22_49 ( .A(u5_mult_82_ab_22__49_), .B(
        u5_mult_82_CARRYB_21__49_), .CI(u5_mult_82_SUMB_21__50_), .CO(
        u5_mult_82_CARRYB_22__49_), .S(u5_mult_82_SUMB_22__49_) );
  FA_X1 u5_mult_82_S2_22_48 ( .A(u5_mult_82_ab_22__48_), .B(
        u5_mult_82_CARRYB_21__48_), .CI(u5_mult_82_SUMB_21__49_), .CO(
        u5_mult_82_CARRYB_22__48_), .S(u5_mult_82_SUMB_22__48_) );
  FA_X1 u5_mult_82_S2_22_47 ( .A(u5_mult_82_ab_22__47_), .B(
        u5_mult_82_CARRYB_21__47_), .CI(u5_mult_82_SUMB_21__48_), .CO(
        u5_mult_82_CARRYB_22__47_), .S(u5_mult_82_SUMB_22__47_) );
  FA_X1 u5_mult_82_S2_22_46 ( .A(u5_mult_82_ab_22__46_), .B(
        u5_mult_82_CARRYB_21__46_), .CI(u5_mult_82_SUMB_21__47_), .CO(
        u5_mult_82_CARRYB_22__46_), .S(u5_mult_82_SUMB_22__46_) );
  FA_X1 u5_mult_82_S2_22_45 ( .A(u5_mult_82_ab_22__45_), .B(
        u5_mult_82_CARRYB_21__45_), .CI(u5_mult_82_SUMB_21__46_), .CO(
        u5_mult_82_CARRYB_22__45_), .S(u5_mult_82_SUMB_22__45_) );
  FA_X1 u5_mult_82_S2_22_44 ( .A(u5_mult_82_ab_22__44_), .B(
        u5_mult_82_CARRYB_21__44_), .CI(u5_mult_82_SUMB_21__45_), .CO(
        u5_mult_82_CARRYB_22__44_), .S(u5_mult_82_SUMB_22__44_) );
  FA_X1 u5_mult_82_S2_22_43 ( .A(u5_mult_82_ab_22__43_), .B(
        u5_mult_82_CARRYB_21__43_), .CI(u5_mult_82_SUMB_21__44_), .CO(
        u5_mult_82_CARRYB_22__43_), .S(u5_mult_82_SUMB_22__43_) );
  FA_X1 u5_mult_82_S2_22_42 ( .A(u5_mult_82_ab_22__42_), .B(
        u5_mult_82_CARRYB_21__42_), .CI(u5_mult_82_SUMB_21__43_), .CO(
        u5_mult_82_CARRYB_22__42_), .S(u5_mult_82_SUMB_22__42_) );
  FA_X1 u5_mult_82_S2_22_41 ( .A(u5_mult_82_ab_22__41_), .B(
        u5_mult_82_CARRYB_21__41_), .CI(u5_mult_82_SUMB_21__42_), .CO(
        u5_mult_82_CARRYB_22__41_), .S(u5_mult_82_SUMB_22__41_) );
  FA_X1 u5_mult_82_S2_22_40 ( .A(u5_mult_82_ab_22__40_), .B(
        u5_mult_82_CARRYB_21__40_), .CI(u5_mult_82_SUMB_21__41_), .CO(
        u5_mult_82_CARRYB_22__40_), .S(u5_mult_82_SUMB_22__40_) );
  FA_X1 u5_mult_82_S2_22_39 ( .A(u5_mult_82_ab_22__39_), .B(
        u5_mult_82_CARRYB_21__39_), .CI(u5_mult_82_SUMB_21__40_), .CO(
        u5_mult_82_CARRYB_22__39_), .S(u5_mult_82_SUMB_22__39_) );
  FA_X1 u5_mult_82_S2_22_38 ( .A(u5_mult_82_ab_22__38_), .B(
        u5_mult_82_CARRYB_21__38_), .CI(u5_mult_82_SUMB_21__39_), .CO(
        u5_mult_82_CARRYB_22__38_), .S(u5_mult_82_SUMB_22__38_) );
  FA_X1 u5_mult_82_S2_22_37 ( .A(u5_mult_82_ab_22__37_), .B(
        u5_mult_82_CARRYB_21__37_), .CI(u5_mult_82_SUMB_21__38_), .CO(
        u5_mult_82_CARRYB_22__37_), .S(u5_mult_82_SUMB_22__37_) );
  FA_X1 u5_mult_82_S2_22_36 ( .A(u5_mult_82_ab_22__36_), .B(
        u5_mult_82_CARRYB_21__36_), .CI(u5_mult_82_SUMB_21__37_), .CO(
        u5_mult_82_CARRYB_22__36_), .S(u5_mult_82_SUMB_22__36_) );
  FA_X1 u5_mult_82_S2_22_35 ( .A(u5_mult_82_ab_22__35_), .B(
        u5_mult_82_CARRYB_21__35_), .CI(u5_mult_82_SUMB_21__36_), .CO(
        u5_mult_82_CARRYB_22__35_), .S(u5_mult_82_SUMB_22__35_) );
  FA_X1 u5_mult_82_S2_22_34 ( .A(u5_mult_82_ab_22__34_), .B(
        u5_mult_82_CARRYB_21__34_), .CI(u5_mult_82_SUMB_21__35_), .CO(
        u5_mult_82_CARRYB_22__34_), .S(u5_mult_82_SUMB_22__34_) );
  FA_X1 u5_mult_82_S2_22_33 ( .A(u5_mult_82_ab_22__33_), .B(
        u5_mult_82_CARRYB_21__33_), .CI(u5_mult_82_SUMB_21__34_), .CO(
        u5_mult_82_CARRYB_22__33_), .S(u5_mult_82_SUMB_22__33_) );
  FA_X1 u5_mult_82_S2_22_32 ( .A(u5_mult_82_ab_22__32_), .B(
        u5_mult_82_CARRYB_21__32_), .CI(u5_mult_82_SUMB_21__33_), .CO(
        u5_mult_82_CARRYB_22__32_), .S(u5_mult_82_SUMB_22__32_) );
  FA_X1 u5_mult_82_S2_22_31 ( .A(u5_mult_82_ab_22__31_), .B(
        u5_mult_82_CARRYB_21__31_), .CI(u5_mult_82_SUMB_21__32_), .CO(
        u5_mult_82_CARRYB_22__31_), .S(u5_mult_82_SUMB_22__31_) );
  FA_X1 u5_mult_82_S2_22_30 ( .A(u5_mult_82_ab_22__30_), .B(
        u5_mult_82_CARRYB_21__30_), .CI(u5_mult_82_SUMB_21__31_), .CO(
        u5_mult_82_CARRYB_22__30_), .S(u5_mult_82_SUMB_22__30_) );
  FA_X1 u5_mult_82_S2_22_29 ( .A(u5_mult_82_ab_22__29_), .B(
        u5_mult_82_CARRYB_21__29_), .CI(u5_mult_82_SUMB_21__30_), .CO(
        u5_mult_82_CARRYB_22__29_), .S(u5_mult_82_SUMB_22__29_) );
  FA_X1 u5_mult_82_S2_22_28 ( .A(u5_mult_82_ab_22__28_), .B(
        u5_mult_82_CARRYB_21__28_), .CI(u5_mult_82_SUMB_21__29_), .CO(
        u5_mult_82_CARRYB_22__28_), .S(u5_mult_82_SUMB_22__28_) );
  FA_X1 u5_mult_82_S2_22_27 ( .A(u5_mult_82_ab_22__27_), .B(
        u5_mult_82_CARRYB_21__27_), .CI(u5_mult_82_SUMB_21__28_), .CO(
        u5_mult_82_CARRYB_22__27_), .S(u5_mult_82_SUMB_22__27_) );
  FA_X1 u5_mult_82_S2_22_26 ( .A(u5_mult_82_ab_22__26_), .B(
        u5_mult_82_CARRYB_21__26_), .CI(u5_mult_82_SUMB_21__27_), .CO(
        u5_mult_82_CARRYB_22__26_), .S(u5_mult_82_SUMB_22__26_) );
  FA_X1 u5_mult_82_S2_22_25 ( .A(u5_mult_82_ab_22__25_), .B(
        u5_mult_82_CARRYB_21__25_), .CI(u5_mult_82_SUMB_21__26_), .CO(
        u5_mult_82_CARRYB_22__25_), .S(u5_mult_82_SUMB_22__25_) );
  FA_X1 u5_mult_82_S2_22_24 ( .A(u5_mult_82_ab_22__24_), .B(
        u5_mult_82_CARRYB_21__24_), .CI(u5_mult_82_SUMB_21__25_), .CO(
        u5_mult_82_CARRYB_22__24_), .S(u5_mult_82_SUMB_22__24_) );
  FA_X1 u5_mult_82_S2_22_23 ( .A(u5_mult_82_ab_22__23_), .B(
        u5_mult_82_CARRYB_21__23_), .CI(u5_mult_82_SUMB_21__24_), .CO(
        u5_mult_82_CARRYB_22__23_), .S(u5_mult_82_SUMB_22__23_) );
  FA_X1 u5_mult_82_S2_22_22 ( .A(u5_mult_82_ab_22__22_), .B(
        u5_mult_82_CARRYB_21__22_), .CI(u5_mult_82_SUMB_21__23_), .CO(
        u5_mult_82_CARRYB_22__22_), .S(u5_mult_82_SUMB_22__22_) );
  FA_X1 u5_mult_82_S2_22_21 ( .A(u5_mult_82_ab_22__21_), .B(
        u5_mult_82_CARRYB_21__21_), .CI(u5_mult_82_SUMB_21__22_), .CO(
        u5_mult_82_CARRYB_22__21_), .S(u5_mult_82_SUMB_22__21_) );
  FA_X1 u5_mult_82_S2_22_20 ( .A(u5_mult_82_ab_22__20_), .B(
        u5_mult_82_CARRYB_21__20_), .CI(u5_mult_82_SUMB_21__21_), .CO(
        u5_mult_82_CARRYB_22__20_), .S(u5_mult_82_SUMB_22__20_) );
  FA_X1 u5_mult_82_S2_22_19 ( .A(u5_mult_82_ab_22__19_), .B(
        u5_mult_82_CARRYB_21__19_), .CI(u5_mult_82_SUMB_21__20_), .CO(
        u5_mult_82_CARRYB_22__19_), .S(u5_mult_82_SUMB_22__19_) );
  FA_X1 u5_mult_82_S2_22_18 ( .A(u5_mult_82_ab_22__18_), .B(
        u5_mult_82_CARRYB_21__18_), .CI(u5_mult_82_SUMB_21__19_), .CO(
        u5_mult_82_CARRYB_22__18_), .S(u5_mult_82_SUMB_22__18_) );
  FA_X1 u5_mult_82_S2_22_17 ( .A(u5_mult_82_ab_22__17_), .B(
        u5_mult_82_CARRYB_21__17_), .CI(u5_mult_82_SUMB_21__18_), .CO(
        u5_mult_82_CARRYB_22__17_), .S(u5_mult_82_SUMB_22__17_) );
  FA_X1 u5_mult_82_S2_22_16 ( .A(u5_mult_82_ab_22__16_), .B(
        u5_mult_82_CARRYB_21__16_), .CI(u5_mult_82_SUMB_21__17_), .CO(
        u5_mult_82_CARRYB_22__16_), .S(u5_mult_82_SUMB_22__16_) );
  FA_X1 u5_mult_82_S2_22_15 ( .A(u5_mult_82_ab_22__15_), .B(
        u5_mult_82_CARRYB_21__15_), .CI(u5_mult_82_SUMB_21__16_), .CO(
        u5_mult_82_CARRYB_22__15_), .S(u5_mult_82_SUMB_22__15_) );
  FA_X1 u5_mult_82_S2_22_14 ( .A(u5_mult_82_ab_22__14_), .B(
        u5_mult_82_CARRYB_21__14_), .CI(u5_mult_82_SUMB_21__15_), .CO(
        u5_mult_82_CARRYB_22__14_), .S(u5_mult_82_SUMB_22__14_) );
  FA_X1 u5_mult_82_S2_22_13 ( .A(u5_mult_82_ab_22__13_), .B(
        u5_mult_82_CARRYB_21__13_), .CI(u5_mult_82_SUMB_21__14_), .CO(
        u5_mult_82_CARRYB_22__13_), .S(u5_mult_82_SUMB_22__13_) );
  FA_X1 u5_mult_82_S2_22_12 ( .A(u5_mult_82_ab_22__12_), .B(
        u5_mult_82_CARRYB_21__12_), .CI(u5_mult_82_SUMB_21__13_), .CO(
        u5_mult_82_CARRYB_22__12_), .S(u5_mult_82_SUMB_22__12_) );
  FA_X1 u5_mult_82_S2_22_11 ( .A(u5_mult_82_ab_22__11_), .B(
        u5_mult_82_CARRYB_21__11_), .CI(u5_mult_82_SUMB_21__12_), .CO(
        u5_mult_82_CARRYB_22__11_), .S(u5_mult_82_SUMB_22__11_) );
  FA_X1 u5_mult_82_S2_22_10 ( .A(u5_mult_82_ab_22__10_), .B(
        u5_mult_82_CARRYB_21__10_), .CI(u5_mult_82_SUMB_21__11_), .CO(
        u5_mult_82_CARRYB_22__10_), .S(u5_mult_82_SUMB_22__10_) );
  FA_X1 u5_mult_82_S2_22_9 ( .A(u5_mult_82_ab_22__9_), .B(
        u5_mult_82_CARRYB_21__9_), .CI(u5_mult_82_SUMB_21__10_), .CO(
        u5_mult_82_CARRYB_22__9_), .S(u5_mult_82_SUMB_22__9_) );
  FA_X1 u5_mult_82_S2_22_8 ( .A(u5_mult_82_ab_22__8_), .B(
        u5_mult_82_CARRYB_21__8_), .CI(u5_mult_82_SUMB_21__9_), .CO(
        u5_mult_82_CARRYB_22__8_), .S(u5_mult_82_SUMB_22__8_) );
  FA_X1 u5_mult_82_S2_22_7 ( .A(u5_mult_82_ab_22__7_), .B(
        u5_mult_82_CARRYB_21__7_), .CI(u5_mult_82_SUMB_21__8_), .CO(
        u5_mult_82_CARRYB_22__7_), .S(u5_mult_82_SUMB_22__7_) );
  FA_X1 u5_mult_82_S2_22_6 ( .A(u5_mult_82_ab_22__6_), .B(
        u5_mult_82_CARRYB_21__6_), .CI(u5_mult_82_SUMB_21__7_), .CO(
        u5_mult_82_CARRYB_22__6_), .S(u5_mult_82_SUMB_22__6_) );
  FA_X1 u5_mult_82_S2_22_5 ( .A(u5_mult_82_ab_22__5_), .B(
        u5_mult_82_CARRYB_21__5_), .CI(u5_mult_82_SUMB_21__6_), .CO(
        u5_mult_82_CARRYB_22__5_), .S(u5_mult_82_SUMB_22__5_) );
  FA_X1 u5_mult_82_S2_22_4 ( .A(u5_mult_82_ab_22__4_), .B(
        u5_mult_82_CARRYB_21__4_), .CI(u5_mult_82_SUMB_21__5_), .CO(
        u5_mult_82_CARRYB_22__4_), .S(u5_mult_82_SUMB_22__4_) );
  FA_X1 u5_mult_82_S2_22_3 ( .A(u5_mult_82_ab_22__3_), .B(
        u5_mult_82_CARRYB_21__3_), .CI(u5_mult_82_SUMB_21__4_), .CO(
        u5_mult_82_CARRYB_22__3_), .S(u5_mult_82_SUMB_22__3_) );
  FA_X1 u5_mult_82_S2_22_2 ( .A(u5_mult_82_ab_22__2_), .B(
        u5_mult_82_CARRYB_21__2_), .CI(u5_mult_82_SUMB_21__3_), .CO(
        u5_mult_82_CARRYB_22__2_), .S(u5_mult_82_SUMB_22__2_) );
  FA_X1 u5_mult_82_S2_22_1 ( .A(u5_mult_82_ab_22__1_), .B(
        u5_mult_82_CARRYB_21__1_), .CI(u5_mult_82_SUMB_21__2_), .CO(
        u5_mult_82_CARRYB_22__1_), .S(u5_mult_82_SUMB_22__1_) );
  FA_X1 u5_mult_82_S1_22_0 ( .A(u5_mult_82_ab_22__0_), .B(
        u5_mult_82_CARRYB_21__0_), .CI(u5_mult_82_SUMB_21__1_), .CO(
        u5_mult_82_CARRYB_22__0_), .S(u5_N22) );
  FA_X1 u5_mult_82_S3_23_51 ( .A(u5_mult_82_ab_23__51_), .B(
        u5_mult_82_CARRYB_22__51_), .CI(u5_mult_82_ab_22__52_), .CO(
        u5_mult_82_CARRYB_23__51_), .S(u5_mult_82_SUMB_23__51_) );
  FA_X1 u5_mult_82_S2_23_50 ( .A(u5_mult_82_ab_23__50_), .B(
        u5_mult_82_CARRYB_22__50_), .CI(u5_mult_82_SUMB_22__51_), .CO(
        u5_mult_82_CARRYB_23__50_), .S(u5_mult_82_SUMB_23__50_) );
  FA_X1 u5_mult_82_S2_23_49 ( .A(u5_mult_82_ab_23__49_), .B(
        u5_mult_82_CARRYB_22__49_), .CI(u5_mult_82_SUMB_22__50_), .CO(
        u5_mult_82_CARRYB_23__49_), .S(u5_mult_82_SUMB_23__49_) );
  FA_X1 u5_mult_82_S2_23_48 ( .A(u5_mult_82_ab_23__48_), .B(
        u5_mult_82_CARRYB_22__48_), .CI(u5_mult_82_SUMB_22__49_), .CO(
        u5_mult_82_CARRYB_23__48_), .S(u5_mult_82_SUMB_23__48_) );
  FA_X1 u5_mult_82_S2_23_47 ( .A(u5_mult_82_ab_23__47_), .B(
        u5_mult_82_CARRYB_22__47_), .CI(u5_mult_82_SUMB_22__48_), .CO(
        u5_mult_82_CARRYB_23__47_), .S(u5_mult_82_SUMB_23__47_) );
  FA_X1 u5_mult_82_S2_23_46 ( .A(u5_mult_82_ab_23__46_), .B(
        u5_mult_82_CARRYB_22__46_), .CI(u5_mult_82_SUMB_22__47_), .CO(
        u5_mult_82_CARRYB_23__46_), .S(u5_mult_82_SUMB_23__46_) );
  FA_X1 u5_mult_82_S2_23_45 ( .A(u5_mult_82_ab_23__45_), .B(
        u5_mult_82_CARRYB_22__45_), .CI(u5_mult_82_SUMB_22__46_), .CO(
        u5_mult_82_CARRYB_23__45_), .S(u5_mult_82_SUMB_23__45_) );
  FA_X1 u5_mult_82_S2_23_44 ( .A(u5_mult_82_ab_23__44_), .B(
        u5_mult_82_CARRYB_22__44_), .CI(u5_mult_82_SUMB_22__45_), .CO(
        u5_mult_82_CARRYB_23__44_), .S(u5_mult_82_SUMB_23__44_) );
  FA_X1 u5_mult_82_S2_23_43 ( .A(u5_mult_82_ab_23__43_), .B(
        u5_mult_82_CARRYB_22__43_), .CI(u5_mult_82_SUMB_22__44_), .CO(
        u5_mult_82_CARRYB_23__43_), .S(u5_mult_82_SUMB_23__43_) );
  FA_X1 u5_mult_82_S2_23_42 ( .A(u5_mult_82_ab_23__42_), .B(
        u5_mult_82_CARRYB_22__42_), .CI(u5_mult_82_SUMB_22__43_), .CO(
        u5_mult_82_CARRYB_23__42_), .S(u5_mult_82_SUMB_23__42_) );
  FA_X1 u5_mult_82_S2_23_41 ( .A(u5_mult_82_ab_23__41_), .B(
        u5_mult_82_CARRYB_22__41_), .CI(u5_mult_82_SUMB_22__42_), .CO(
        u5_mult_82_CARRYB_23__41_), .S(u5_mult_82_SUMB_23__41_) );
  FA_X1 u5_mult_82_S2_23_40 ( .A(u5_mult_82_ab_23__40_), .B(
        u5_mult_82_CARRYB_22__40_), .CI(u5_mult_82_SUMB_22__41_), .CO(
        u5_mult_82_CARRYB_23__40_), .S(u5_mult_82_SUMB_23__40_) );
  FA_X1 u5_mult_82_S2_23_39 ( .A(u5_mult_82_ab_23__39_), .B(
        u5_mult_82_CARRYB_22__39_), .CI(u5_mult_82_SUMB_22__40_), .CO(
        u5_mult_82_CARRYB_23__39_), .S(u5_mult_82_SUMB_23__39_) );
  FA_X1 u5_mult_82_S2_23_38 ( .A(u5_mult_82_ab_23__38_), .B(
        u5_mult_82_CARRYB_22__38_), .CI(u5_mult_82_SUMB_22__39_), .CO(
        u5_mult_82_CARRYB_23__38_), .S(u5_mult_82_SUMB_23__38_) );
  FA_X1 u5_mult_82_S2_23_37 ( .A(u5_mult_82_ab_23__37_), .B(
        u5_mult_82_CARRYB_22__37_), .CI(u5_mult_82_SUMB_22__38_), .CO(
        u5_mult_82_CARRYB_23__37_), .S(u5_mult_82_SUMB_23__37_) );
  FA_X1 u5_mult_82_S2_23_36 ( .A(u5_mult_82_ab_23__36_), .B(
        u5_mult_82_CARRYB_22__36_), .CI(u5_mult_82_SUMB_22__37_), .CO(
        u5_mult_82_CARRYB_23__36_), .S(u5_mult_82_SUMB_23__36_) );
  FA_X1 u5_mult_82_S2_23_35 ( .A(u5_mult_82_ab_23__35_), .B(
        u5_mult_82_CARRYB_22__35_), .CI(u5_mult_82_SUMB_22__36_), .CO(
        u5_mult_82_CARRYB_23__35_), .S(u5_mult_82_SUMB_23__35_) );
  FA_X1 u5_mult_82_S2_23_34 ( .A(u5_mult_82_ab_23__34_), .B(
        u5_mult_82_CARRYB_22__34_), .CI(u5_mult_82_SUMB_22__35_), .CO(
        u5_mult_82_CARRYB_23__34_), .S(u5_mult_82_SUMB_23__34_) );
  FA_X1 u5_mult_82_S2_23_33 ( .A(u5_mult_82_ab_23__33_), .B(
        u5_mult_82_CARRYB_22__33_), .CI(u5_mult_82_SUMB_22__34_), .CO(
        u5_mult_82_CARRYB_23__33_), .S(u5_mult_82_SUMB_23__33_) );
  FA_X1 u5_mult_82_S2_23_32 ( .A(u5_mult_82_ab_23__32_), .B(
        u5_mult_82_CARRYB_22__32_), .CI(u5_mult_82_SUMB_22__33_), .CO(
        u5_mult_82_CARRYB_23__32_), .S(u5_mult_82_SUMB_23__32_) );
  FA_X1 u5_mult_82_S2_23_31 ( .A(u5_mult_82_ab_23__31_), .B(
        u5_mult_82_CARRYB_22__31_), .CI(u5_mult_82_SUMB_22__32_), .CO(
        u5_mult_82_CARRYB_23__31_), .S(u5_mult_82_SUMB_23__31_) );
  FA_X1 u5_mult_82_S2_23_30 ( .A(u5_mult_82_ab_23__30_), .B(
        u5_mult_82_CARRYB_22__30_), .CI(u5_mult_82_SUMB_22__31_), .CO(
        u5_mult_82_CARRYB_23__30_), .S(u5_mult_82_SUMB_23__30_) );
  FA_X1 u5_mult_82_S2_23_29 ( .A(u5_mult_82_ab_23__29_), .B(
        u5_mult_82_CARRYB_22__29_), .CI(u5_mult_82_SUMB_22__30_), .CO(
        u5_mult_82_CARRYB_23__29_), .S(u5_mult_82_SUMB_23__29_) );
  FA_X1 u5_mult_82_S2_23_28 ( .A(u5_mult_82_ab_23__28_), .B(
        u5_mult_82_CARRYB_22__28_), .CI(u5_mult_82_SUMB_22__29_), .CO(
        u5_mult_82_CARRYB_23__28_), .S(u5_mult_82_SUMB_23__28_) );
  FA_X1 u5_mult_82_S2_23_27 ( .A(u5_mult_82_ab_23__27_), .B(
        u5_mult_82_CARRYB_22__27_), .CI(u5_mult_82_SUMB_22__28_), .CO(
        u5_mult_82_CARRYB_23__27_), .S(u5_mult_82_SUMB_23__27_) );
  FA_X1 u5_mult_82_S2_23_26 ( .A(u5_mult_82_ab_23__26_), .B(
        u5_mult_82_CARRYB_22__26_), .CI(u5_mult_82_SUMB_22__27_), .CO(
        u5_mult_82_CARRYB_23__26_), .S(u5_mult_82_SUMB_23__26_) );
  FA_X1 u5_mult_82_S2_23_25 ( .A(u5_mult_82_ab_23__25_), .B(
        u5_mult_82_CARRYB_22__25_), .CI(u5_mult_82_SUMB_22__26_), .CO(
        u5_mult_82_CARRYB_23__25_), .S(u5_mult_82_SUMB_23__25_) );
  FA_X1 u5_mult_82_S2_23_24 ( .A(u5_mult_82_ab_23__24_), .B(
        u5_mult_82_CARRYB_22__24_), .CI(u5_mult_82_SUMB_22__25_), .CO(
        u5_mult_82_CARRYB_23__24_), .S(u5_mult_82_SUMB_23__24_) );
  FA_X1 u5_mult_82_S2_23_23 ( .A(u5_mult_82_ab_23__23_), .B(
        u5_mult_82_CARRYB_22__23_), .CI(u5_mult_82_SUMB_22__24_), .CO(
        u5_mult_82_CARRYB_23__23_), .S(u5_mult_82_SUMB_23__23_) );
  FA_X1 u5_mult_82_S2_23_22 ( .A(u5_mult_82_ab_23__22_), .B(
        u5_mult_82_CARRYB_22__22_), .CI(u5_mult_82_SUMB_22__23_), .CO(
        u5_mult_82_CARRYB_23__22_), .S(u5_mult_82_SUMB_23__22_) );
  FA_X1 u5_mult_82_S2_23_21 ( .A(u5_mult_82_ab_23__21_), .B(
        u5_mult_82_CARRYB_22__21_), .CI(u5_mult_82_SUMB_22__22_), .CO(
        u5_mult_82_CARRYB_23__21_), .S(u5_mult_82_SUMB_23__21_) );
  FA_X1 u5_mult_82_S2_23_20 ( .A(u5_mult_82_ab_23__20_), .B(
        u5_mult_82_CARRYB_22__20_), .CI(u5_mult_82_SUMB_22__21_), .CO(
        u5_mult_82_CARRYB_23__20_), .S(u5_mult_82_SUMB_23__20_) );
  FA_X1 u5_mult_82_S2_23_19 ( .A(u5_mult_82_ab_23__19_), .B(
        u5_mult_82_CARRYB_22__19_), .CI(u5_mult_82_SUMB_22__20_), .CO(
        u5_mult_82_CARRYB_23__19_), .S(u5_mult_82_SUMB_23__19_) );
  FA_X1 u5_mult_82_S2_23_18 ( .A(u5_mult_82_ab_23__18_), .B(
        u5_mult_82_CARRYB_22__18_), .CI(u5_mult_82_SUMB_22__19_), .CO(
        u5_mult_82_CARRYB_23__18_), .S(u5_mult_82_SUMB_23__18_) );
  FA_X1 u5_mult_82_S2_23_17 ( .A(u5_mult_82_ab_23__17_), .B(
        u5_mult_82_CARRYB_22__17_), .CI(u5_mult_82_SUMB_22__18_), .CO(
        u5_mult_82_CARRYB_23__17_), .S(u5_mult_82_SUMB_23__17_) );
  FA_X1 u5_mult_82_S2_23_16 ( .A(u5_mult_82_ab_23__16_), .B(
        u5_mult_82_CARRYB_22__16_), .CI(u5_mult_82_SUMB_22__17_), .CO(
        u5_mult_82_CARRYB_23__16_), .S(u5_mult_82_SUMB_23__16_) );
  FA_X1 u5_mult_82_S2_23_15 ( .A(u5_mult_82_ab_23__15_), .B(
        u5_mult_82_CARRYB_22__15_), .CI(u5_mult_82_SUMB_22__16_), .CO(
        u5_mult_82_CARRYB_23__15_), .S(u5_mult_82_SUMB_23__15_) );
  FA_X1 u5_mult_82_S2_23_14 ( .A(u5_mult_82_ab_23__14_), .B(
        u5_mult_82_CARRYB_22__14_), .CI(u5_mult_82_SUMB_22__15_), .CO(
        u5_mult_82_CARRYB_23__14_), .S(u5_mult_82_SUMB_23__14_) );
  FA_X1 u5_mult_82_S2_23_13 ( .A(u5_mult_82_ab_23__13_), .B(
        u5_mult_82_CARRYB_22__13_), .CI(u5_mult_82_SUMB_22__14_), .CO(
        u5_mult_82_CARRYB_23__13_), .S(u5_mult_82_SUMB_23__13_) );
  FA_X1 u5_mult_82_S2_23_12 ( .A(u5_mult_82_ab_23__12_), .B(
        u5_mult_82_CARRYB_22__12_), .CI(u5_mult_82_SUMB_22__13_), .CO(
        u5_mult_82_CARRYB_23__12_), .S(u5_mult_82_SUMB_23__12_) );
  FA_X1 u5_mult_82_S2_23_11 ( .A(u5_mult_82_ab_23__11_), .B(
        u5_mult_82_CARRYB_22__11_), .CI(u5_mult_82_SUMB_22__12_), .CO(
        u5_mult_82_CARRYB_23__11_), .S(u5_mult_82_SUMB_23__11_) );
  FA_X1 u5_mult_82_S2_23_10 ( .A(u5_mult_82_ab_23__10_), .B(
        u5_mult_82_CARRYB_22__10_), .CI(u5_mult_82_SUMB_22__11_), .CO(
        u5_mult_82_CARRYB_23__10_), .S(u5_mult_82_SUMB_23__10_) );
  FA_X1 u5_mult_82_S2_23_9 ( .A(u5_mult_82_ab_23__9_), .B(
        u5_mult_82_CARRYB_22__9_), .CI(u5_mult_82_SUMB_22__10_), .CO(
        u5_mult_82_CARRYB_23__9_), .S(u5_mult_82_SUMB_23__9_) );
  FA_X1 u5_mult_82_S2_23_8 ( .A(u5_mult_82_ab_23__8_), .B(
        u5_mult_82_CARRYB_22__8_), .CI(u5_mult_82_SUMB_22__9_), .CO(
        u5_mult_82_CARRYB_23__8_), .S(u5_mult_82_SUMB_23__8_) );
  FA_X1 u5_mult_82_S2_23_7 ( .A(u5_mult_82_ab_23__7_), .B(
        u5_mult_82_CARRYB_22__7_), .CI(u5_mult_82_SUMB_22__8_), .CO(
        u5_mult_82_CARRYB_23__7_), .S(u5_mult_82_SUMB_23__7_) );
  FA_X1 u5_mult_82_S2_23_6 ( .A(u5_mult_82_ab_23__6_), .B(
        u5_mult_82_CARRYB_22__6_), .CI(u5_mult_82_SUMB_22__7_), .CO(
        u5_mult_82_CARRYB_23__6_), .S(u5_mult_82_SUMB_23__6_) );
  FA_X1 u5_mult_82_S2_23_5 ( .A(u5_mult_82_ab_23__5_), .B(
        u5_mult_82_CARRYB_22__5_), .CI(u5_mult_82_SUMB_22__6_), .CO(
        u5_mult_82_CARRYB_23__5_), .S(u5_mult_82_SUMB_23__5_) );
  FA_X1 u5_mult_82_S2_23_4 ( .A(u5_mult_82_ab_23__4_), .B(
        u5_mult_82_CARRYB_22__4_), .CI(u5_mult_82_SUMB_22__5_), .CO(
        u5_mult_82_CARRYB_23__4_), .S(u5_mult_82_SUMB_23__4_) );
  FA_X1 u5_mult_82_S2_23_3 ( .A(u5_mult_82_ab_23__3_), .B(
        u5_mult_82_CARRYB_22__3_), .CI(u5_mult_82_SUMB_22__4_), .CO(
        u5_mult_82_CARRYB_23__3_), .S(u5_mult_82_SUMB_23__3_) );
  FA_X1 u5_mult_82_S2_23_2 ( .A(u5_mult_82_ab_23__2_), .B(
        u5_mult_82_CARRYB_22__2_), .CI(u5_mult_82_SUMB_22__3_), .CO(
        u5_mult_82_CARRYB_23__2_), .S(u5_mult_82_SUMB_23__2_) );
  FA_X1 u5_mult_82_S2_23_1 ( .A(u5_mult_82_ab_23__1_), .B(
        u5_mult_82_CARRYB_22__1_), .CI(u5_mult_82_SUMB_22__2_), .CO(
        u5_mult_82_CARRYB_23__1_), .S(u5_mult_82_SUMB_23__1_) );
  FA_X1 u5_mult_82_S1_23_0 ( .A(u5_mult_82_ab_23__0_), .B(
        u5_mult_82_CARRYB_22__0_), .CI(u5_mult_82_SUMB_22__1_), .CO(
        u5_mult_82_CARRYB_23__0_), .S(u5_N23) );
  FA_X1 u5_mult_82_S3_24_51 ( .A(u5_mult_82_ab_24__51_), .B(
        u5_mult_82_CARRYB_23__51_), .CI(u5_mult_82_ab_23__52_), .CO(
        u5_mult_82_CARRYB_24__51_), .S(u5_mult_82_SUMB_24__51_) );
  FA_X1 u5_mult_82_S2_24_50 ( .A(u5_mult_82_ab_24__50_), .B(
        u5_mult_82_CARRYB_23__50_), .CI(u5_mult_82_SUMB_23__51_), .CO(
        u5_mult_82_CARRYB_24__50_), .S(u5_mult_82_SUMB_24__50_) );
  FA_X1 u5_mult_82_S2_24_49 ( .A(u5_mult_82_ab_24__49_), .B(
        u5_mult_82_CARRYB_23__49_), .CI(u5_mult_82_SUMB_23__50_), .CO(
        u5_mult_82_CARRYB_24__49_), .S(u5_mult_82_SUMB_24__49_) );
  FA_X1 u5_mult_82_S2_24_48 ( .A(u5_mult_82_ab_24__48_), .B(
        u5_mult_82_CARRYB_23__48_), .CI(u5_mult_82_SUMB_23__49_), .CO(
        u5_mult_82_CARRYB_24__48_), .S(u5_mult_82_SUMB_24__48_) );
  FA_X1 u5_mult_82_S2_24_47 ( .A(u5_mult_82_ab_24__47_), .B(
        u5_mult_82_CARRYB_23__47_), .CI(u5_mult_82_SUMB_23__48_), .CO(
        u5_mult_82_CARRYB_24__47_), .S(u5_mult_82_SUMB_24__47_) );
  FA_X1 u5_mult_82_S2_24_46 ( .A(u5_mult_82_ab_24__46_), .B(
        u5_mult_82_CARRYB_23__46_), .CI(u5_mult_82_SUMB_23__47_), .CO(
        u5_mult_82_CARRYB_24__46_), .S(u5_mult_82_SUMB_24__46_) );
  FA_X1 u5_mult_82_S2_24_45 ( .A(u5_mult_82_ab_24__45_), .B(
        u5_mult_82_CARRYB_23__45_), .CI(u5_mult_82_SUMB_23__46_), .CO(
        u5_mult_82_CARRYB_24__45_), .S(u5_mult_82_SUMB_24__45_) );
  FA_X1 u5_mult_82_S2_24_44 ( .A(u5_mult_82_ab_24__44_), .B(
        u5_mult_82_CARRYB_23__44_), .CI(u5_mult_82_SUMB_23__45_), .CO(
        u5_mult_82_CARRYB_24__44_), .S(u5_mult_82_SUMB_24__44_) );
  FA_X1 u5_mult_82_S2_24_43 ( .A(u5_mult_82_ab_24__43_), .B(
        u5_mult_82_CARRYB_23__43_), .CI(u5_mult_82_SUMB_23__44_), .CO(
        u5_mult_82_CARRYB_24__43_), .S(u5_mult_82_SUMB_24__43_) );
  FA_X1 u5_mult_82_S2_24_42 ( .A(u5_mult_82_ab_24__42_), .B(
        u5_mult_82_CARRYB_23__42_), .CI(u5_mult_82_SUMB_23__43_), .CO(
        u5_mult_82_CARRYB_24__42_), .S(u5_mult_82_SUMB_24__42_) );
  FA_X1 u5_mult_82_S2_24_41 ( .A(u5_mult_82_ab_24__41_), .B(
        u5_mult_82_CARRYB_23__41_), .CI(u5_mult_82_SUMB_23__42_), .CO(
        u5_mult_82_CARRYB_24__41_), .S(u5_mult_82_SUMB_24__41_) );
  FA_X1 u5_mult_82_S2_24_40 ( .A(u5_mult_82_ab_24__40_), .B(
        u5_mult_82_CARRYB_23__40_), .CI(u5_mult_82_SUMB_23__41_), .CO(
        u5_mult_82_CARRYB_24__40_), .S(u5_mult_82_SUMB_24__40_) );
  FA_X1 u5_mult_82_S2_24_39 ( .A(u5_mult_82_ab_24__39_), .B(
        u5_mult_82_CARRYB_23__39_), .CI(u5_mult_82_SUMB_23__40_), .CO(
        u5_mult_82_CARRYB_24__39_), .S(u5_mult_82_SUMB_24__39_) );
  FA_X1 u5_mult_82_S2_24_38 ( .A(u5_mult_82_ab_24__38_), .B(
        u5_mult_82_CARRYB_23__38_), .CI(u5_mult_82_SUMB_23__39_), .CO(
        u5_mult_82_CARRYB_24__38_), .S(u5_mult_82_SUMB_24__38_) );
  FA_X1 u5_mult_82_S2_24_37 ( .A(u5_mult_82_ab_24__37_), .B(
        u5_mult_82_CARRYB_23__37_), .CI(u5_mult_82_SUMB_23__38_), .CO(
        u5_mult_82_CARRYB_24__37_), .S(u5_mult_82_SUMB_24__37_) );
  FA_X1 u5_mult_82_S2_24_36 ( .A(u5_mult_82_ab_24__36_), .B(
        u5_mult_82_CARRYB_23__36_), .CI(u5_mult_82_SUMB_23__37_), .CO(
        u5_mult_82_CARRYB_24__36_), .S(u5_mult_82_SUMB_24__36_) );
  FA_X1 u5_mult_82_S2_24_35 ( .A(u5_mult_82_ab_24__35_), .B(
        u5_mult_82_CARRYB_23__35_), .CI(u5_mult_82_SUMB_23__36_), .CO(
        u5_mult_82_CARRYB_24__35_), .S(u5_mult_82_SUMB_24__35_) );
  FA_X1 u5_mult_82_S2_24_34 ( .A(u5_mult_82_ab_24__34_), .B(
        u5_mult_82_CARRYB_23__34_), .CI(u5_mult_82_SUMB_23__35_), .CO(
        u5_mult_82_CARRYB_24__34_), .S(u5_mult_82_SUMB_24__34_) );
  FA_X1 u5_mult_82_S2_24_33 ( .A(u5_mult_82_ab_24__33_), .B(
        u5_mult_82_CARRYB_23__33_), .CI(u5_mult_82_SUMB_23__34_), .CO(
        u5_mult_82_CARRYB_24__33_), .S(u5_mult_82_SUMB_24__33_) );
  FA_X1 u5_mult_82_S2_24_32 ( .A(u5_mult_82_ab_24__32_), .B(
        u5_mult_82_CARRYB_23__32_), .CI(u5_mult_82_SUMB_23__33_), .CO(
        u5_mult_82_CARRYB_24__32_), .S(u5_mult_82_SUMB_24__32_) );
  FA_X1 u5_mult_82_S2_24_31 ( .A(u5_mult_82_ab_24__31_), .B(
        u5_mult_82_CARRYB_23__31_), .CI(u5_mult_82_SUMB_23__32_), .CO(
        u5_mult_82_CARRYB_24__31_), .S(u5_mult_82_SUMB_24__31_) );
  FA_X1 u5_mult_82_S2_24_30 ( .A(u5_mult_82_ab_24__30_), .B(
        u5_mult_82_CARRYB_23__30_), .CI(u5_mult_82_SUMB_23__31_), .CO(
        u5_mult_82_CARRYB_24__30_), .S(u5_mult_82_SUMB_24__30_) );
  FA_X1 u5_mult_82_S2_24_29 ( .A(u5_mult_82_ab_24__29_), .B(
        u5_mult_82_CARRYB_23__29_), .CI(u5_mult_82_SUMB_23__30_), .CO(
        u5_mult_82_CARRYB_24__29_), .S(u5_mult_82_SUMB_24__29_) );
  FA_X1 u5_mult_82_S2_24_28 ( .A(u5_mult_82_ab_24__28_), .B(
        u5_mult_82_CARRYB_23__28_), .CI(u5_mult_82_SUMB_23__29_), .CO(
        u5_mult_82_CARRYB_24__28_), .S(u5_mult_82_SUMB_24__28_) );
  FA_X1 u5_mult_82_S2_24_27 ( .A(u5_mult_82_ab_24__27_), .B(
        u5_mult_82_CARRYB_23__27_), .CI(u5_mult_82_SUMB_23__28_), .CO(
        u5_mult_82_CARRYB_24__27_), .S(u5_mult_82_SUMB_24__27_) );
  FA_X1 u5_mult_82_S2_24_26 ( .A(u5_mult_82_ab_24__26_), .B(
        u5_mult_82_CARRYB_23__26_), .CI(u5_mult_82_SUMB_23__27_), .CO(
        u5_mult_82_CARRYB_24__26_), .S(u5_mult_82_SUMB_24__26_) );
  FA_X1 u5_mult_82_S2_24_25 ( .A(u5_mult_82_ab_24__25_), .B(
        u5_mult_82_CARRYB_23__25_), .CI(u5_mult_82_SUMB_23__26_), .CO(
        u5_mult_82_CARRYB_24__25_), .S(u5_mult_82_SUMB_24__25_) );
  FA_X1 u5_mult_82_S2_24_24 ( .A(u5_mult_82_ab_24__24_), .B(
        u5_mult_82_CARRYB_23__24_), .CI(u5_mult_82_SUMB_23__25_), .CO(
        u5_mult_82_CARRYB_24__24_), .S(u5_mult_82_SUMB_24__24_) );
  FA_X1 u5_mult_82_S2_24_23 ( .A(u5_mult_82_ab_24__23_), .B(
        u5_mult_82_CARRYB_23__23_), .CI(u5_mult_82_SUMB_23__24_), .CO(
        u5_mult_82_CARRYB_24__23_), .S(u5_mult_82_SUMB_24__23_) );
  FA_X1 u5_mult_82_S2_24_22 ( .A(u5_mult_82_ab_24__22_), .B(
        u5_mult_82_CARRYB_23__22_), .CI(u5_mult_82_SUMB_23__23_), .CO(
        u5_mult_82_CARRYB_24__22_), .S(u5_mult_82_SUMB_24__22_) );
  FA_X1 u5_mult_82_S2_24_21 ( .A(u5_mult_82_ab_24__21_), .B(
        u5_mult_82_CARRYB_23__21_), .CI(u5_mult_82_SUMB_23__22_), .CO(
        u5_mult_82_CARRYB_24__21_), .S(u5_mult_82_SUMB_24__21_) );
  FA_X1 u5_mult_82_S2_24_20 ( .A(u5_mult_82_ab_24__20_), .B(
        u5_mult_82_CARRYB_23__20_), .CI(u5_mult_82_SUMB_23__21_), .CO(
        u5_mult_82_CARRYB_24__20_), .S(u5_mult_82_SUMB_24__20_) );
  FA_X1 u5_mult_82_S2_24_19 ( .A(u5_mult_82_ab_24__19_), .B(
        u5_mult_82_CARRYB_23__19_), .CI(u5_mult_82_SUMB_23__20_), .CO(
        u5_mult_82_CARRYB_24__19_), .S(u5_mult_82_SUMB_24__19_) );
  FA_X1 u5_mult_82_S2_24_18 ( .A(u5_mult_82_ab_24__18_), .B(
        u5_mult_82_CARRYB_23__18_), .CI(u5_mult_82_SUMB_23__19_), .CO(
        u5_mult_82_CARRYB_24__18_), .S(u5_mult_82_SUMB_24__18_) );
  FA_X1 u5_mult_82_S2_24_17 ( .A(u5_mult_82_ab_24__17_), .B(
        u5_mult_82_CARRYB_23__17_), .CI(u5_mult_82_SUMB_23__18_), .CO(
        u5_mult_82_CARRYB_24__17_), .S(u5_mult_82_SUMB_24__17_) );
  FA_X1 u5_mult_82_S2_24_16 ( .A(u5_mult_82_ab_24__16_), .B(
        u5_mult_82_CARRYB_23__16_), .CI(u5_mult_82_SUMB_23__17_), .CO(
        u5_mult_82_CARRYB_24__16_), .S(u5_mult_82_SUMB_24__16_) );
  FA_X1 u5_mult_82_S2_24_15 ( .A(u5_mult_82_ab_24__15_), .B(
        u5_mult_82_CARRYB_23__15_), .CI(u5_mult_82_SUMB_23__16_), .CO(
        u5_mult_82_CARRYB_24__15_), .S(u5_mult_82_SUMB_24__15_) );
  FA_X1 u5_mult_82_S2_24_14 ( .A(u5_mult_82_ab_24__14_), .B(
        u5_mult_82_CARRYB_23__14_), .CI(u5_mult_82_SUMB_23__15_), .CO(
        u5_mult_82_CARRYB_24__14_), .S(u5_mult_82_SUMB_24__14_) );
  FA_X1 u5_mult_82_S2_24_13 ( .A(u5_mult_82_ab_24__13_), .B(
        u5_mult_82_CARRYB_23__13_), .CI(u5_mult_82_SUMB_23__14_), .CO(
        u5_mult_82_CARRYB_24__13_), .S(u5_mult_82_SUMB_24__13_) );
  FA_X1 u5_mult_82_S2_24_12 ( .A(u5_mult_82_ab_24__12_), .B(
        u5_mult_82_CARRYB_23__12_), .CI(u5_mult_82_SUMB_23__13_), .CO(
        u5_mult_82_CARRYB_24__12_), .S(u5_mult_82_SUMB_24__12_) );
  FA_X1 u5_mult_82_S2_24_11 ( .A(u5_mult_82_ab_24__11_), .B(
        u5_mult_82_CARRYB_23__11_), .CI(u5_mult_82_SUMB_23__12_), .CO(
        u5_mult_82_CARRYB_24__11_), .S(u5_mult_82_SUMB_24__11_) );
  FA_X1 u5_mult_82_S2_24_10 ( .A(u5_mult_82_ab_24__10_), .B(
        u5_mult_82_CARRYB_23__10_), .CI(u5_mult_82_SUMB_23__11_), .CO(
        u5_mult_82_CARRYB_24__10_), .S(u5_mult_82_SUMB_24__10_) );
  FA_X1 u5_mult_82_S2_24_9 ( .A(u5_mult_82_ab_24__9_), .B(
        u5_mult_82_CARRYB_23__9_), .CI(u5_mult_82_SUMB_23__10_), .CO(
        u5_mult_82_CARRYB_24__9_), .S(u5_mult_82_SUMB_24__9_) );
  FA_X1 u5_mult_82_S2_24_8 ( .A(u5_mult_82_ab_24__8_), .B(
        u5_mult_82_CARRYB_23__8_), .CI(u5_mult_82_SUMB_23__9_), .CO(
        u5_mult_82_CARRYB_24__8_), .S(u5_mult_82_SUMB_24__8_) );
  FA_X1 u5_mult_82_S2_24_7 ( .A(u5_mult_82_ab_24__7_), .B(
        u5_mult_82_CARRYB_23__7_), .CI(u5_mult_82_SUMB_23__8_), .CO(
        u5_mult_82_CARRYB_24__7_), .S(u5_mult_82_SUMB_24__7_) );
  FA_X1 u5_mult_82_S2_24_6 ( .A(u5_mult_82_ab_24__6_), .B(
        u5_mult_82_CARRYB_23__6_), .CI(u5_mult_82_SUMB_23__7_), .CO(
        u5_mult_82_CARRYB_24__6_), .S(u5_mult_82_SUMB_24__6_) );
  FA_X1 u5_mult_82_S2_24_5 ( .A(u5_mult_82_ab_24__5_), .B(
        u5_mult_82_CARRYB_23__5_), .CI(u5_mult_82_SUMB_23__6_), .CO(
        u5_mult_82_CARRYB_24__5_), .S(u5_mult_82_SUMB_24__5_) );
  FA_X1 u5_mult_82_S2_24_4 ( .A(u5_mult_82_ab_24__4_), .B(
        u5_mult_82_CARRYB_23__4_), .CI(u5_mult_82_SUMB_23__5_), .CO(
        u5_mult_82_CARRYB_24__4_), .S(u5_mult_82_SUMB_24__4_) );
  FA_X1 u5_mult_82_S2_24_3 ( .A(u5_mult_82_ab_24__3_), .B(
        u5_mult_82_CARRYB_23__3_), .CI(u5_mult_82_SUMB_23__4_), .CO(
        u5_mult_82_CARRYB_24__3_), .S(u5_mult_82_SUMB_24__3_) );
  FA_X1 u5_mult_82_S2_24_2 ( .A(u5_mult_82_ab_24__2_), .B(
        u5_mult_82_CARRYB_23__2_), .CI(u5_mult_82_SUMB_23__3_), .CO(
        u5_mult_82_CARRYB_24__2_), .S(u5_mult_82_SUMB_24__2_) );
  FA_X1 u5_mult_82_S2_24_1 ( .A(u5_mult_82_ab_24__1_), .B(
        u5_mult_82_CARRYB_23__1_), .CI(u5_mult_82_SUMB_23__2_), .CO(
        u5_mult_82_CARRYB_24__1_), .S(u5_mult_82_SUMB_24__1_) );
  FA_X1 u5_mult_82_S1_24_0 ( .A(u5_mult_82_ab_24__0_), .B(
        u5_mult_82_CARRYB_23__0_), .CI(u5_mult_82_SUMB_23__1_), .CO(
        u5_mult_82_CARRYB_24__0_), .S(u5_N24) );
  FA_X1 u5_mult_82_S3_25_51 ( .A(u5_mult_82_ab_25__51_), .B(
        u5_mult_82_CARRYB_24__51_), .CI(u5_mult_82_ab_24__52_), .CO(
        u5_mult_82_CARRYB_25__51_), .S(u5_mult_82_SUMB_25__51_) );
  FA_X1 u5_mult_82_S2_25_50 ( .A(u5_mult_82_ab_25__50_), .B(
        u5_mult_82_CARRYB_24__50_), .CI(u5_mult_82_SUMB_24__51_), .CO(
        u5_mult_82_CARRYB_25__50_), .S(u5_mult_82_SUMB_25__50_) );
  FA_X1 u5_mult_82_S2_25_49 ( .A(u5_mult_82_ab_25__49_), .B(
        u5_mult_82_CARRYB_24__49_), .CI(u5_mult_82_SUMB_24__50_), .CO(
        u5_mult_82_CARRYB_25__49_), .S(u5_mult_82_SUMB_25__49_) );
  FA_X1 u5_mult_82_S2_25_48 ( .A(u5_mult_82_ab_25__48_), .B(
        u5_mult_82_CARRYB_24__48_), .CI(u5_mult_82_SUMB_24__49_), .CO(
        u5_mult_82_CARRYB_25__48_), .S(u5_mult_82_SUMB_25__48_) );
  FA_X1 u5_mult_82_S2_25_47 ( .A(u5_mult_82_ab_25__47_), .B(
        u5_mult_82_CARRYB_24__47_), .CI(u5_mult_82_SUMB_24__48_), .CO(
        u5_mult_82_CARRYB_25__47_), .S(u5_mult_82_SUMB_25__47_) );
  FA_X1 u5_mult_82_S2_25_46 ( .A(u5_mult_82_ab_25__46_), .B(
        u5_mult_82_CARRYB_24__46_), .CI(u5_mult_82_SUMB_24__47_), .CO(
        u5_mult_82_CARRYB_25__46_), .S(u5_mult_82_SUMB_25__46_) );
  FA_X1 u5_mult_82_S2_25_45 ( .A(u5_mult_82_ab_25__45_), .B(
        u5_mult_82_CARRYB_24__45_), .CI(u5_mult_82_SUMB_24__46_), .CO(
        u5_mult_82_CARRYB_25__45_), .S(u5_mult_82_SUMB_25__45_) );
  FA_X1 u5_mult_82_S2_25_44 ( .A(u5_mult_82_ab_25__44_), .B(
        u5_mult_82_CARRYB_24__44_), .CI(u5_mult_82_SUMB_24__45_), .CO(
        u5_mult_82_CARRYB_25__44_), .S(u5_mult_82_SUMB_25__44_) );
  FA_X1 u5_mult_82_S2_25_43 ( .A(u5_mult_82_ab_25__43_), .B(
        u5_mult_82_CARRYB_24__43_), .CI(u5_mult_82_SUMB_24__44_), .CO(
        u5_mult_82_CARRYB_25__43_), .S(u5_mult_82_SUMB_25__43_) );
  FA_X1 u5_mult_82_S2_25_42 ( .A(u5_mult_82_ab_25__42_), .B(
        u5_mult_82_CARRYB_24__42_), .CI(u5_mult_82_SUMB_24__43_), .CO(
        u5_mult_82_CARRYB_25__42_), .S(u5_mult_82_SUMB_25__42_) );
  FA_X1 u5_mult_82_S2_25_41 ( .A(u5_mult_82_ab_25__41_), .B(
        u5_mult_82_CARRYB_24__41_), .CI(u5_mult_82_SUMB_24__42_), .CO(
        u5_mult_82_CARRYB_25__41_), .S(u5_mult_82_SUMB_25__41_) );
  FA_X1 u5_mult_82_S2_25_40 ( .A(u5_mult_82_ab_25__40_), .B(
        u5_mult_82_CARRYB_24__40_), .CI(u5_mult_82_SUMB_24__41_), .CO(
        u5_mult_82_CARRYB_25__40_), .S(u5_mult_82_SUMB_25__40_) );
  FA_X1 u5_mult_82_S2_25_39 ( .A(u5_mult_82_ab_25__39_), .B(
        u5_mult_82_CARRYB_24__39_), .CI(u5_mult_82_SUMB_24__40_), .CO(
        u5_mult_82_CARRYB_25__39_), .S(u5_mult_82_SUMB_25__39_) );
  FA_X1 u5_mult_82_S2_25_38 ( .A(u5_mult_82_ab_25__38_), .B(
        u5_mult_82_CARRYB_24__38_), .CI(u5_mult_82_SUMB_24__39_), .CO(
        u5_mult_82_CARRYB_25__38_), .S(u5_mult_82_SUMB_25__38_) );
  FA_X1 u5_mult_82_S2_25_37 ( .A(u5_mult_82_ab_25__37_), .B(
        u5_mult_82_CARRYB_24__37_), .CI(u5_mult_82_SUMB_24__38_), .CO(
        u5_mult_82_CARRYB_25__37_), .S(u5_mult_82_SUMB_25__37_) );
  FA_X1 u5_mult_82_S2_25_36 ( .A(u5_mult_82_ab_25__36_), .B(
        u5_mult_82_CARRYB_24__36_), .CI(u5_mult_82_SUMB_24__37_), .CO(
        u5_mult_82_CARRYB_25__36_), .S(u5_mult_82_SUMB_25__36_) );
  FA_X1 u5_mult_82_S2_25_35 ( .A(u5_mult_82_ab_25__35_), .B(
        u5_mult_82_CARRYB_24__35_), .CI(u5_mult_82_SUMB_24__36_), .CO(
        u5_mult_82_CARRYB_25__35_), .S(u5_mult_82_SUMB_25__35_) );
  FA_X1 u5_mult_82_S2_25_34 ( .A(u5_mult_82_ab_25__34_), .B(
        u5_mult_82_CARRYB_24__34_), .CI(u5_mult_82_SUMB_24__35_), .CO(
        u5_mult_82_CARRYB_25__34_), .S(u5_mult_82_SUMB_25__34_) );
  FA_X1 u5_mult_82_S2_25_33 ( .A(u5_mult_82_ab_25__33_), .B(
        u5_mult_82_CARRYB_24__33_), .CI(u5_mult_82_SUMB_24__34_), .CO(
        u5_mult_82_CARRYB_25__33_), .S(u5_mult_82_SUMB_25__33_) );
  FA_X1 u5_mult_82_S2_25_32 ( .A(u5_mult_82_ab_25__32_), .B(
        u5_mult_82_CARRYB_24__32_), .CI(u5_mult_82_SUMB_24__33_), .CO(
        u5_mult_82_CARRYB_25__32_), .S(u5_mult_82_SUMB_25__32_) );
  FA_X1 u5_mult_82_S2_25_31 ( .A(u5_mult_82_ab_25__31_), .B(
        u5_mult_82_CARRYB_24__31_), .CI(u5_mult_82_SUMB_24__32_), .CO(
        u5_mult_82_CARRYB_25__31_), .S(u5_mult_82_SUMB_25__31_) );
  FA_X1 u5_mult_82_S2_25_30 ( .A(u5_mult_82_ab_25__30_), .B(
        u5_mult_82_CARRYB_24__30_), .CI(u5_mult_82_SUMB_24__31_), .CO(
        u5_mult_82_CARRYB_25__30_), .S(u5_mult_82_SUMB_25__30_) );
  FA_X1 u5_mult_82_S2_25_29 ( .A(u5_mult_82_ab_25__29_), .B(
        u5_mult_82_CARRYB_24__29_), .CI(u5_mult_82_SUMB_24__30_), .CO(
        u5_mult_82_CARRYB_25__29_), .S(u5_mult_82_SUMB_25__29_) );
  FA_X1 u5_mult_82_S2_25_28 ( .A(u5_mult_82_ab_25__28_), .B(
        u5_mult_82_CARRYB_24__28_), .CI(u5_mult_82_SUMB_24__29_), .CO(
        u5_mult_82_CARRYB_25__28_), .S(u5_mult_82_SUMB_25__28_) );
  FA_X1 u5_mult_82_S2_25_27 ( .A(u5_mult_82_ab_25__27_), .B(
        u5_mult_82_CARRYB_24__27_), .CI(u5_mult_82_SUMB_24__28_), .CO(
        u5_mult_82_CARRYB_25__27_), .S(u5_mult_82_SUMB_25__27_) );
  FA_X1 u5_mult_82_S2_25_26 ( .A(u5_mult_82_ab_25__26_), .B(
        u5_mult_82_CARRYB_24__26_), .CI(u5_mult_82_SUMB_24__27_), .CO(
        u5_mult_82_CARRYB_25__26_), .S(u5_mult_82_SUMB_25__26_) );
  FA_X1 u5_mult_82_S2_25_25 ( .A(u5_mult_82_ab_25__25_), .B(
        u5_mult_82_CARRYB_24__25_), .CI(u5_mult_82_SUMB_24__26_), .CO(
        u5_mult_82_CARRYB_25__25_), .S(u5_mult_82_SUMB_25__25_) );
  FA_X1 u5_mult_82_S2_25_24 ( .A(u5_mult_82_ab_25__24_), .B(
        u5_mult_82_CARRYB_24__24_), .CI(u5_mult_82_SUMB_24__25_), .CO(
        u5_mult_82_CARRYB_25__24_), .S(u5_mult_82_SUMB_25__24_) );
  FA_X1 u5_mult_82_S2_25_23 ( .A(u5_mult_82_ab_25__23_), .B(
        u5_mult_82_CARRYB_24__23_), .CI(u5_mult_82_SUMB_24__24_), .CO(
        u5_mult_82_CARRYB_25__23_), .S(u5_mult_82_SUMB_25__23_) );
  FA_X1 u5_mult_82_S2_25_22 ( .A(u5_mult_82_ab_25__22_), .B(
        u5_mult_82_CARRYB_24__22_), .CI(u5_mult_82_SUMB_24__23_), .CO(
        u5_mult_82_CARRYB_25__22_), .S(u5_mult_82_SUMB_25__22_) );
  FA_X1 u5_mult_82_S2_25_21 ( .A(u5_mult_82_ab_25__21_), .B(
        u5_mult_82_CARRYB_24__21_), .CI(u5_mult_82_SUMB_24__22_), .CO(
        u5_mult_82_CARRYB_25__21_), .S(u5_mult_82_SUMB_25__21_) );
  FA_X1 u5_mult_82_S2_25_20 ( .A(u5_mult_82_ab_25__20_), .B(
        u5_mult_82_CARRYB_24__20_), .CI(u5_mult_82_SUMB_24__21_), .CO(
        u5_mult_82_CARRYB_25__20_), .S(u5_mult_82_SUMB_25__20_) );
  FA_X1 u5_mult_82_S2_25_19 ( .A(u5_mult_82_ab_25__19_), .B(
        u5_mult_82_CARRYB_24__19_), .CI(u5_mult_82_SUMB_24__20_), .CO(
        u5_mult_82_CARRYB_25__19_), .S(u5_mult_82_SUMB_25__19_) );
  FA_X1 u5_mult_82_S2_25_18 ( .A(u5_mult_82_ab_25__18_), .B(
        u5_mult_82_CARRYB_24__18_), .CI(u5_mult_82_SUMB_24__19_), .CO(
        u5_mult_82_CARRYB_25__18_), .S(u5_mult_82_SUMB_25__18_) );
  FA_X1 u5_mult_82_S2_25_17 ( .A(u5_mult_82_ab_25__17_), .B(
        u5_mult_82_CARRYB_24__17_), .CI(u5_mult_82_SUMB_24__18_), .CO(
        u5_mult_82_CARRYB_25__17_), .S(u5_mult_82_SUMB_25__17_) );
  FA_X1 u5_mult_82_S2_25_16 ( .A(u5_mult_82_ab_25__16_), .B(
        u5_mult_82_CARRYB_24__16_), .CI(u5_mult_82_SUMB_24__17_), .CO(
        u5_mult_82_CARRYB_25__16_), .S(u5_mult_82_SUMB_25__16_) );
  FA_X1 u5_mult_82_S2_25_15 ( .A(u5_mult_82_ab_25__15_), .B(
        u5_mult_82_CARRYB_24__15_), .CI(u5_mult_82_SUMB_24__16_), .CO(
        u5_mult_82_CARRYB_25__15_), .S(u5_mult_82_SUMB_25__15_) );
  FA_X1 u5_mult_82_S2_25_14 ( .A(u5_mult_82_ab_25__14_), .B(
        u5_mult_82_CARRYB_24__14_), .CI(u5_mult_82_SUMB_24__15_), .CO(
        u5_mult_82_CARRYB_25__14_), .S(u5_mult_82_SUMB_25__14_) );
  FA_X1 u5_mult_82_S2_25_13 ( .A(u5_mult_82_ab_25__13_), .B(
        u5_mult_82_CARRYB_24__13_), .CI(u5_mult_82_SUMB_24__14_), .CO(
        u5_mult_82_CARRYB_25__13_), .S(u5_mult_82_SUMB_25__13_) );
  FA_X1 u5_mult_82_S2_25_12 ( .A(u5_mult_82_ab_25__12_), .B(
        u5_mult_82_CARRYB_24__12_), .CI(u5_mult_82_SUMB_24__13_), .CO(
        u5_mult_82_CARRYB_25__12_), .S(u5_mult_82_SUMB_25__12_) );
  FA_X1 u5_mult_82_S2_25_11 ( .A(u5_mult_82_ab_25__11_), .B(
        u5_mult_82_CARRYB_24__11_), .CI(u5_mult_82_SUMB_24__12_), .CO(
        u5_mult_82_CARRYB_25__11_), .S(u5_mult_82_SUMB_25__11_) );
  FA_X1 u5_mult_82_S2_25_10 ( .A(u5_mult_82_ab_25__10_), .B(
        u5_mult_82_CARRYB_24__10_), .CI(u5_mult_82_SUMB_24__11_), .CO(
        u5_mult_82_CARRYB_25__10_), .S(u5_mult_82_SUMB_25__10_) );
  FA_X1 u5_mult_82_S2_25_9 ( .A(u5_mult_82_ab_25__9_), .B(
        u5_mult_82_CARRYB_24__9_), .CI(u5_mult_82_SUMB_24__10_), .CO(
        u5_mult_82_CARRYB_25__9_), .S(u5_mult_82_SUMB_25__9_) );
  FA_X1 u5_mult_82_S2_25_8 ( .A(u5_mult_82_ab_25__8_), .B(
        u5_mult_82_CARRYB_24__8_), .CI(u5_mult_82_SUMB_24__9_), .CO(
        u5_mult_82_CARRYB_25__8_), .S(u5_mult_82_SUMB_25__8_) );
  FA_X1 u5_mult_82_S2_25_7 ( .A(u5_mult_82_ab_25__7_), .B(
        u5_mult_82_CARRYB_24__7_), .CI(u5_mult_82_SUMB_24__8_), .CO(
        u5_mult_82_CARRYB_25__7_), .S(u5_mult_82_SUMB_25__7_) );
  FA_X1 u5_mult_82_S2_25_6 ( .A(u5_mult_82_ab_25__6_), .B(
        u5_mult_82_CARRYB_24__6_), .CI(u5_mult_82_SUMB_24__7_), .CO(
        u5_mult_82_CARRYB_25__6_), .S(u5_mult_82_SUMB_25__6_) );
  FA_X1 u5_mult_82_S2_25_5 ( .A(u5_mult_82_ab_25__5_), .B(
        u5_mult_82_CARRYB_24__5_), .CI(u5_mult_82_SUMB_24__6_), .CO(
        u5_mult_82_CARRYB_25__5_), .S(u5_mult_82_SUMB_25__5_) );
  FA_X1 u5_mult_82_S2_25_4 ( .A(u5_mult_82_ab_25__4_), .B(
        u5_mult_82_CARRYB_24__4_), .CI(u5_mult_82_SUMB_24__5_), .CO(
        u5_mult_82_CARRYB_25__4_), .S(u5_mult_82_SUMB_25__4_) );
  FA_X1 u5_mult_82_S2_25_3 ( .A(u5_mult_82_ab_25__3_), .B(
        u5_mult_82_CARRYB_24__3_), .CI(u5_mult_82_SUMB_24__4_), .CO(
        u5_mult_82_CARRYB_25__3_), .S(u5_mult_82_SUMB_25__3_) );
  FA_X1 u5_mult_82_S2_25_2 ( .A(u5_mult_82_ab_25__2_), .B(
        u5_mult_82_CARRYB_24__2_), .CI(u5_mult_82_SUMB_24__3_), .CO(
        u5_mult_82_CARRYB_25__2_), .S(u5_mult_82_SUMB_25__2_) );
  FA_X1 u5_mult_82_S2_25_1 ( .A(u5_mult_82_ab_25__1_), .B(
        u5_mult_82_CARRYB_24__1_), .CI(u5_mult_82_SUMB_24__2_), .CO(
        u5_mult_82_CARRYB_25__1_), .S(u5_mult_82_SUMB_25__1_) );
  FA_X1 u5_mult_82_S1_25_0 ( .A(u5_mult_82_ab_25__0_), .B(
        u5_mult_82_CARRYB_24__0_), .CI(u5_mult_82_SUMB_24__1_), .CO(
        u5_mult_82_CARRYB_25__0_), .S(u5_N25) );
  FA_X1 u5_mult_82_S3_26_51 ( .A(u5_mult_82_ab_26__51_), .B(
        u5_mult_82_CARRYB_25__51_), .CI(u5_mult_82_ab_25__52_), .CO(
        u5_mult_82_CARRYB_26__51_), .S(u5_mult_82_SUMB_26__51_) );
  FA_X1 u5_mult_82_S2_26_50 ( .A(u5_mult_82_ab_26__50_), .B(
        u5_mult_82_CARRYB_25__50_), .CI(u5_mult_82_SUMB_25__51_), .CO(
        u5_mult_82_CARRYB_26__50_), .S(u5_mult_82_SUMB_26__50_) );
  FA_X1 u5_mult_82_S2_26_49 ( .A(u5_mult_82_ab_26__49_), .B(
        u5_mult_82_CARRYB_25__49_), .CI(u5_mult_82_SUMB_25__50_), .CO(
        u5_mult_82_CARRYB_26__49_), .S(u5_mult_82_SUMB_26__49_) );
  FA_X1 u5_mult_82_S2_26_48 ( .A(u5_mult_82_ab_26__48_), .B(
        u5_mult_82_CARRYB_25__48_), .CI(u5_mult_82_SUMB_25__49_), .CO(
        u5_mult_82_CARRYB_26__48_), .S(u5_mult_82_SUMB_26__48_) );
  FA_X1 u5_mult_82_S2_26_47 ( .A(u5_mult_82_ab_26__47_), .B(
        u5_mult_82_CARRYB_25__47_), .CI(u5_mult_82_SUMB_25__48_), .CO(
        u5_mult_82_CARRYB_26__47_), .S(u5_mult_82_SUMB_26__47_) );
  FA_X1 u5_mult_82_S2_26_46 ( .A(u5_mult_82_ab_26__46_), .B(
        u5_mult_82_CARRYB_25__46_), .CI(u5_mult_82_SUMB_25__47_), .CO(
        u5_mult_82_CARRYB_26__46_), .S(u5_mult_82_SUMB_26__46_) );
  FA_X1 u5_mult_82_S2_26_45 ( .A(u5_mult_82_ab_26__45_), .B(
        u5_mult_82_CARRYB_25__45_), .CI(u5_mult_82_SUMB_25__46_), .CO(
        u5_mult_82_CARRYB_26__45_), .S(u5_mult_82_SUMB_26__45_) );
  FA_X1 u5_mult_82_S2_26_44 ( .A(u5_mult_82_ab_26__44_), .B(
        u5_mult_82_CARRYB_25__44_), .CI(u5_mult_82_SUMB_25__45_), .CO(
        u5_mult_82_CARRYB_26__44_), .S(u5_mult_82_SUMB_26__44_) );
  FA_X1 u5_mult_82_S2_26_43 ( .A(u5_mult_82_ab_26__43_), .B(
        u5_mult_82_CARRYB_25__43_), .CI(u5_mult_82_SUMB_25__44_), .CO(
        u5_mult_82_CARRYB_26__43_), .S(u5_mult_82_SUMB_26__43_) );
  FA_X1 u5_mult_82_S2_26_42 ( .A(u5_mult_82_ab_26__42_), .B(
        u5_mult_82_CARRYB_25__42_), .CI(u5_mult_82_SUMB_25__43_), .CO(
        u5_mult_82_CARRYB_26__42_), .S(u5_mult_82_SUMB_26__42_) );
  FA_X1 u5_mult_82_S2_26_41 ( .A(u5_mult_82_ab_26__41_), .B(
        u5_mult_82_CARRYB_25__41_), .CI(u5_mult_82_SUMB_25__42_), .CO(
        u5_mult_82_CARRYB_26__41_), .S(u5_mult_82_SUMB_26__41_) );
  FA_X1 u5_mult_82_S2_26_40 ( .A(u5_mult_82_ab_26__40_), .B(
        u5_mult_82_CARRYB_25__40_), .CI(u5_mult_82_SUMB_25__41_), .CO(
        u5_mult_82_CARRYB_26__40_), .S(u5_mult_82_SUMB_26__40_) );
  FA_X1 u5_mult_82_S2_26_39 ( .A(u5_mult_82_ab_26__39_), .B(
        u5_mult_82_CARRYB_25__39_), .CI(u5_mult_82_SUMB_25__40_), .CO(
        u5_mult_82_CARRYB_26__39_), .S(u5_mult_82_SUMB_26__39_) );
  FA_X1 u5_mult_82_S2_26_38 ( .A(u5_mult_82_ab_26__38_), .B(
        u5_mult_82_CARRYB_25__38_), .CI(u5_mult_82_SUMB_25__39_), .CO(
        u5_mult_82_CARRYB_26__38_), .S(u5_mult_82_SUMB_26__38_) );
  FA_X1 u5_mult_82_S2_26_37 ( .A(u5_mult_82_ab_26__37_), .B(
        u5_mult_82_CARRYB_25__37_), .CI(u5_mult_82_SUMB_25__38_), .CO(
        u5_mult_82_CARRYB_26__37_), .S(u5_mult_82_SUMB_26__37_) );
  FA_X1 u5_mult_82_S2_26_36 ( .A(u5_mult_82_ab_26__36_), .B(
        u5_mult_82_CARRYB_25__36_), .CI(u5_mult_82_SUMB_25__37_), .CO(
        u5_mult_82_CARRYB_26__36_), .S(u5_mult_82_SUMB_26__36_) );
  FA_X1 u5_mult_82_S2_26_35 ( .A(u5_mult_82_ab_26__35_), .B(
        u5_mult_82_CARRYB_25__35_), .CI(u5_mult_82_SUMB_25__36_), .CO(
        u5_mult_82_CARRYB_26__35_), .S(u5_mult_82_SUMB_26__35_) );
  FA_X1 u5_mult_82_S2_26_34 ( .A(u5_mult_82_ab_26__34_), .B(
        u5_mult_82_CARRYB_25__34_), .CI(u5_mult_82_SUMB_25__35_), .CO(
        u5_mult_82_CARRYB_26__34_), .S(u5_mult_82_SUMB_26__34_) );
  FA_X1 u5_mult_82_S2_26_33 ( .A(u5_mult_82_ab_26__33_), .B(
        u5_mult_82_CARRYB_25__33_), .CI(u5_mult_82_SUMB_25__34_), .CO(
        u5_mult_82_CARRYB_26__33_), .S(u5_mult_82_SUMB_26__33_) );
  FA_X1 u5_mult_82_S2_26_32 ( .A(u5_mult_82_ab_26__32_), .B(
        u5_mult_82_CARRYB_25__32_), .CI(u5_mult_82_SUMB_25__33_), .CO(
        u5_mult_82_CARRYB_26__32_), .S(u5_mult_82_SUMB_26__32_) );
  FA_X1 u5_mult_82_S2_26_31 ( .A(u5_mult_82_ab_26__31_), .B(
        u5_mult_82_CARRYB_25__31_), .CI(u5_mult_82_SUMB_25__32_), .CO(
        u5_mult_82_CARRYB_26__31_), .S(u5_mult_82_SUMB_26__31_) );
  FA_X1 u5_mult_82_S2_26_30 ( .A(u5_mult_82_ab_26__30_), .B(
        u5_mult_82_CARRYB_25__30_), .CI(u5_mult_82_SUMB_25__31_), .CO(
        u5_mult_82_CARRYB_26__30_), .S(u5_mult_82_SUMB_26__30_) );
  FA_X1 u5_mult_82_S2_26_29 ( .A(u5_mult_82_ab_26__29_), .B(
        u5_mult_82_CARRYB_25__29_), .CI(u5_mult_82_SUMB_25__30_), .CO(
        u5_mult_82_CARRYB_26__29_), .S(u5_mult_82_SUMB_26__29_) );
  FA_X1 u5_mult_82_S2_26_28 ( .A(u5_mult_82_ab_26__28_), .B(
        u5_mult_82_CARRYB_25__28_), .CI(u5_mult_82_SUMB_25__29_), .CO(
        u5_mult_82_CARRYB_26__28_), .S(u5_mult_82_SUMB_26__28_) );
  FA_X1 u5_mult_82_S2_26_27 ( .A(u5_mult_82_ab_26__27_), .B(
        u5_mult_82_CARRYB_25__27_), .CI(u5_mult_82_SUMB_25__28_), .CO(
        u5_mult_82_CARRYB_26__27_), .S(u5_mult_82_SUMB_26__27_) );
  FA_X1 u5_mult_82_S2_26_26 ( .A(u5_mult_82_ab_26__26_), .B(
        u5_mult_82_CARRYB_25__26_), .CI(u5_mult_82_SUMB_25__27_), .CO(
        u5_mult_82_CARRYB_26__26_), .S(u5_mult_82_SUMB_26__26_) );
  FA_X1 u5_mult_82_S2_26_25 ( .A(u5_mult_82_ab_26__25_), .B(
        u5_mult_82_CARRYB_25__25_), .CI(u5_mult_82_SUMB_25__26_), .CO(
        u5_mult_82_CARRYB_26__25_), .S(u5_mult_82_SUMB_26__25_) );
  FA_X1 u5_mult_82_S2_26_24 ( .A(u5_mult_82_ab_26__24_), .B(
        u5_mult_82_CARRYB_25__24_), .CI(u5_mult_82_SUMB_25__25_), .CO(
        u5_mult_82_CARRYB_26__24_), .S(u5_mult_82_SUMB_26__24_) );
  FA_X1 u5_mult_82_S2_26_23 ( .A(u5_mult_82_ab_26__23_), .B(
        u5_mult_82_CARRYB_25__23_), .CI(u5_mult_82_SUMB_25__24_), .CO(
        u5_mult_82_CARRYB_26__23_), .S(u5_mult_82_SUMB_26__23_) );
  FA_X1 u5_mult_82_S2_26_22 ( .A(u5_mult_82_ab_26__22_), .B(
        u5_mult_82_CARRYB_25__22_), .CI(u5_mult_82_SUMB_25__23_), .CO(
        u5_mult_82_CARRYB_26__22_), .S(u5_mult_82_SUMB_26__22_) );
  FA_X1 u5_mult_82_S2_26_21 ( .A(u5_mult_82_ab_26__21_), .B(
        u5_mult_82_CARRYB_25__21_), .CI(u5_mult_82_SUMB_25__22_), .CO(
        u5_mult_82_CARRYB_26__21_), .S(u5_mult_82_SUMB_26__21_) );
  FA_X1 u5_mult_82_S2_26_20 ( .A(u5_mult_82_ab_26__20_), .B(
        u5_mult_82_CARRYB_25__20_), .CI(u5_mult_82_SUMB_25__21_), .CO(
        u5_mult_82_CARRYB_26__20_), .S(u5_mult_82_SUMB_26__20_) );
  FA_X1 u5_mult_82_S2_26_19 ( .A(u5_mult_82_ab_26__19_), .B(
        u5_mult_82_CARRYB_25__19_), .CI(u5_mult_82_SUMB_25__20_), .CO(
        u5_mult_82_CARRYB_26__19_), .S(u5_mult_82_SUMB_26__19_) );
  FA_X1 u5_mult_82_S2_26_18 ( .A(u5_mult_82_ab_26__18_), .B(
        u5_mult_82_CARRYB_25__18_), .CI(u5_mult_82_SUMB_25__19_), .CO(
        u5_mult_82_CARRYB_26__18_), .S(u5_mult_82_SUMB_26__18_) );
  FA_X1 u5_mult_82_S2_26_17 ( .A(u5_mult_82_ab_26__17_), .B(
        u5_mult_82_CARRYB_25__17_), .CI(u5_mult_82_SUMB_25__18_), .CO(
        u5_mult_82_CARRYB_26__17_), .S(u5_mult_82_SUMB_26__17_) );
  FA_X1 u5_mult_82_S2_26_16 ( .A(u5_mult_82_ab_26__16_), .B(
        u5_mult_82_CARRYB_25__16_), .CI(u5_mult_82_SUMB_25__17_), .CO(
        u5_mult_82_CARRYB_26__16_), .S(u5_mult_82_SUMB_26__16_) );
  FA_X1 u5_mult_82_S2_26_15 ( .A(u5_mult_82_ab_26__15_), .B(
        u5_mult_82_CARRYB_25__15_), .CI(u5_mult_82_SUMB_25__16_), .CO(
        u5_mult_82_CARRYB_26__15_), .S(u5_mult_82_SUMB_26__15_) );
  FA_X1 u5_mult_82_S2_26_14 ( .A(u5_mult_82_ab_26__14_), .B(
        u5_mult_82_CARRYB_25__14_), .CI(u5_mult_82_SUMB_25__15_), .CO(
        u5_mult_82_CARRYB_26__14_), .S(u5_mult_82_SUMB_26__14_) );
  FA_X1 u5_mult_82_S2_26_13 ( .A(u5_mult_82_ab_26__13_), .B(
        u5_mult_82_CARRYB_25__13_), .CI(u5_mult_82_SUMB_25__14_), .CO(
        u5_mult_82_CARRYB_26__13_), .S(u5_mult_82_SUMB_26__13_) );
  FA_X1 u5_mult_82_S2_26_12 ( .A(u5_mult_82_ab_26__12_), .B(
        u5_mult_82_CARRYB_25__12_), .CI(u5_mult_82_SUMB_25__13_), .CO(
        u5_mult_82_CARRYB_26__12_), .S(u5_mult_82_SUMB_26__12_) );
  FA_X1 u5_mult_82_S2_26_11 ( .A(u5_mult_82_ab_26__11_), .B(
        u5_mult_82_CARRYB_25__11_), .CI(u5_mult_82_SUMB_25__12_), .CO(
        u5_mult_82_CARRYB_26__11_), .S(u5_mult_82_SUMB_26__11_) );
  FA_X1 u5_mult_82_S2_26_10 ( .A(u5_mult_82_ab_26__10_), .B(
        u5_mult_82_CARRYB_25__10_), .CI(u5_mult_82_SUMB_25__11_), .CO(
        u5_mult_82_CARRYB_26__10_), .S(u5_mult_82_SUMB_26__10_) );
  FA_X1 u5_mult_82_S2_26_9 ( .A(u5_mult_82_ab_26__9_), .B(
        u5_mult_82_CARRYB_25__9_), .CI(u5_mult_82_SUMB_25__10_), .CO(
        u5_mult_82_CARRYB_26__9_), .S(u5_mult_82_SUMB_26__9_) );
  FA_X1 u5_mult_82_S2_26_8 ( .A(u5_mult_82_ab_26__8_), .B(
        u5_mult_82_CARRYB_25__8_), .CI(u5_mult_82_SUMB_25__9_), .CO(
        u5_mult_82_CARRYB_26__8_), .S(u5_mult_82_SUMB_26__8_) );
  FA_X1 u5_mult_82_S2_26_7 ( .A(u5_mult_82_ab_26__7_), .B(
        u5_mult_82_CARRYB_25__7_), .CI(u5_mult_82_SUMB_25__8_), .CO(
        u5_mult_82_CARRYB_26__7_), .S(u5_mult_82_SUMB_26__7_) );
  FA_X1 u5_mult_82_S2_26_6 ( .A(u5_mult_82_ab_26__6_), .B(
        u5_mult_82_CARRYB_25__6_), .CI(u5_mult_82_SUMB_25__7_), .CO(
        u5_mult_82_CARRYB_26__6_), .S(u5_mult_82_SUMB_26__6_) );
  FA_X1 u5_mult_82_S2_26_5 ( .A(u5_mult_82_ab_26__5_), .B(
        u5_mult_82_CARRYB_25__5_), .CI(u5_mult_82_SUMB_25__6_), .CO(
        u5_mult_82_CARRYB_26__5_), .S(u5_mult_82_SUMB_26__5_) );
  FA_X1 u5_mult_82_S2_26_4 ( .A(u5_mult_82_ab_26__4_), .B(
        u5_mult_82_CARRYB_25__4_), .CI(u5_mult_82_SUMB_25__5_), .CO(
        u5_mult_82_CARRYB_26__4_), .S(u5_mult_82_SUMB_26__4_) );
  FA_X1 u5_mult_82_S2_26_3 ( .A(u5_mult_82_ab_26__3_), .B(
        u5_mult_82_CARRYB_25__3_), .CI(u5_mult_82_SUMB_25__4_), .CO(
        u5_mult_82_CARRYB_26__3_), .S(u5_mult_82_SUMB_26__3_) );
  FA_X1 u5_mult_82_S2_26_2 ( .A(u5_mult_82_ab_26__2_), .B(
        u5_mult_82_CARRYB_25__2_), .CI(u5_mult_82_SUMB_25__3_), .CO(
        u5_mult_82_CARRYB_26__2_), .S(u5_mult_82_SUMB_26__2_) );
  FA_X1 u5_mult_82_S2_26_1 ( .A(u5_mult_82_ab_26__1_), .B(
        u5_mult_82_CARRYB_25__1_), .CI(u5_mult_82_SUMB_25__2_), .CO(
        u5_mult_82_CARRYB_26__1_), .S(u5_mult_82_SUMB_26__1_) );
  FA_X1 u5_mult_82_S1_26_0 ( .A(u5_mult_82_ab_26__0_), .B(
        u5_mult_82_CARRYB_25__0_), .CI(u5_mult_82_SUMB_25__1_), .CO(
        u5_mult_82_CARRYB_26__0_), .S(u5_N26) );
  FA_X1 u5_mult_82_S3_27_51 ( .A(u5_mult_82_ab_27__51_), .B(
        u5_mult_82_CARRYB_26__51_), .CI(u5_mult_82_ab_26__52_), .CO(
        u5_mult_82_CARRYB_27__51_), .S(u5_mult_82_SUMB_27__51_) );
  FA_X1 u5_mult_82_S2_27_50 ( .A(u5_mult_82_ab_27__50_), .B(
        u5_mult_82_CARRYB_26__50_), .CI(u5_mult_82_SUMB_26__51_), .CO(
        u5_mult_82_CARRYB_27__50_), .S(u5_mult_82_SUMB_27__50_) );
  FA_X1 u5_mult_82_S2_27_49 ( .A(u5_mult_82_ab_27__49_), .B(
        u5_mult_82_CARRYB_26__49_), .CI(u5_mult_82_SUMB_26__50_), .CO(
        u5_mult_82_CARRYB_27__49_), .S(u5_mult_82_SUMB_27__49_) );
  FA_X1 u5_mult_82_S2_27_48 ( .A(u5_mult_82_ab_27__48_), .B(
        u5_mult_82_CARRYB_26__48_), .CI(u5_mult_82_SUMB_26__49_), .CO(
        u5_mult_82_CARRYB_27__48_), .S(u5_mult_82_SUMB_27__48_) );
  FA_X1 u5_mult_82_S2_27_47 ( .A(u5_mult_82_ab_27__47_), .B(
        u5_mult_82_CARRYB_26__47_), .CI(u5_mult_82_SUMB_26__48_), .CO(
        u5_mult_82_CARRYB_27__47_), .S(u5_mult_82_SUMB_27__47_) );
  FA_X1 u5_mult_82_S2_27_46 ( .A(u5_mult_82_ab_27__46_), .B(
        u5_mult_82_CARRYB_26__46_), .CI(u5_mult_82_SUMB_26__47_), .CO(
        u5_mult_82_CARRYB_27__46_), .S(u5_mult_82_SUMB_27__46_) );
  FA_X1 u5_mult_82_S2_27_45 ( .A(u5_mult_82_ab_27__45_), .B(
        u5_mult_82_CARRYB_26__45_), .CI(u5_mult_82_SUMB_26__46_), .CO(
        u5_mult_82_CARRYB_27__45_), .S(u5_mult_82_SUMB_27__45_) );
  FA_X1 u5_mult_82_S2_27_44 ( .A(u5_mult_82_ab_27__44_), .B(
        u5_mult_82_CARRYB_26__44_), .CI(u5_mult_82_SUMB_26__45_), .CO(
        u5_mult_82_CARRYB_27__44_), .S(u5_mult_82_SUMB_27__44_) );
  FA_X1 u5_mult_82_S2_27_43 ( .A(u5_mult_82_ab_27__43_), .B(
        u5_mult_82_CARRYB_26__43_), .CI(u5_mult_82_SUMB_26__44_), .CO(
        u5_mult_82_CARRYB_27__43_), .S(u5_mult_82_SUMB_27__43_) );
  FA_X1 u5_mult_82_S2_27_42 ( .A(u5_mult_82_ab_27__42_), .B(
        u5_mult_82_CARRYB_26__42_), .CI(u5_mult_82_SUMB_26__43_), .CO(
        u5_mult_82_CARRYB_27__42_), .S(u5_mult_82_SUMB_27__42_) );
  FA_X1 u5_mult_82_S2_27_41 ( .A(u5_mult_82_ab_27__41_), .B(
        u5_mult_82_CARRYB_26__41_), .CI(u5_mult_82_SUMB_26__42_), .CO(
        u5_mult_82_CARRYB_27__41_), .S(u5_mult_82_SUMB_27__41_) );
  FA_X1 u5_mult_82_S2_27_40 ( .A(u5_mult_82_ab_27__40_), .B(
        u5_mult_82_CARRYB_26__40_), .CI(u5_mult_82_SUMB_26__41_), .CO(
        u5_mult_82_CARRYB_27__40_), .S(u5_mult_82_SUMB_27__40_) );
  FA_X1 u5_mult_82_S2_27_39 ( .A(u5_mult_82_ab_27__39_), .B(
        u5_mult_82_CARRYB_26__39_), .CI(u5_mult_82_SUMB_26__40_), .CO(
        u5_mult_82_CARRYB_27__39_), .S(u5_mult_82_SUMB_27__39_) );
  FA_X1 u5_mult_82_S2_27_38 ( .A(u5_mult_82_ab_27__38_), .B(
        u5_mult_82_CARRYB_26__38_), .CI(u5_mult_82_SUMB_26__39_), .CO(
        u5_mult_82_CARRYB_27__38_), .S(u5_mult_82_SUMB_27__38_) );
  FA_X1 u5_mult_82_S2_27_37 ( .A(u5_mult_82_ab_27__37_), .B(
        u5_mult_82_CARRYB_26__37_), .CI(u5_mult_82_SUMB_26__38_), .CO(
        u5_mult_82_CARRYB_27__37_), .S(u5_mult_82_SUMB_27__37_) );
  FA_X1 u5_mult_82_S2_27_36 ( .A(u5_mult_82_ab_27__36_), .B(
        u5_mult_82_CARRYB_26__36_), .CI(u5_mult_82_SUMB_26__37_), .CO(
        u5_mult_82_CARRYB_27__36_), .S(u5_mult_82_SUMB_27__36_) );
  FA_X1 u5_mult_82_S2_27_35 ( .A(u5_mult_82_ab_27__35_), .B(
        u5_mult_82_CARRYB_26__35_), .CI(u5_mult_82_SUMB_26__36_), .CO(
        u5_mult_82_CARRYB_27__35_), .S(u5_mult_82_SUMB_27__35_) );
  FA_X1 u5_mult_82_S2_27_34 ( .A(u5_mult_82_ab_27__34_), .B(
        u5_mult_82_CARRYB_26__34_), .CI(u5_mult_82_SUMB_26__35_), .CO(
        u5_mult_82_CARRYB_27__34_), .S(u5_mult_82_SUMB_27__34_) );
  FA_X1 u5_mult_82_S2_27_33 ( .A(u5_mult_82_ab_27__33_), .B(
        u5_mult_82_CARRYB_26__33_), .CI(u5_mult_82_SUMB_26__34_), .CO(
        u5_mult_82_CARRYB_27__33_), .S(u5_mult_82_SUMB_27__33_) );
  FA_X1 u5_mult_82_S2_27_32 ( .A(u5_mult_82_ab_27__32_), .B(
        u5_mult_82_CARRYB_26__32_), .CI(u5_mult_82_SUMB_26__33_), .CO(
        u5_mult_82_CARRYB_27__32_), .S(u5_mult_82_SUMB_27__32_) );
  FA_X1 u5_mult_82_S2_27_31 ( .A(u5_mult_82_ab_27__31_), .B(
        u5_mult_82_CARRYB_26__31_), .CI(u5_mult_82_SUMB_26__32_), .CO(
        u5_mult_82_CARRYB_27__31_), .S(u5_mult_82_SUMB_27__31_) );
  FA_X1 u5_mult_82_S2_27_30 ( .A(u5_mult_82_ab_27__30_), .B(
        u5_mult_82_CARRYB_26__30_), .CI(u5_mult_82_SUMB_26__31_), .CO(
        u5_mult_82_CARRYB_27__30_), .S(u5_mult_82_SUMB_27__30_) );
  FA_X1 u5_mult_82_S2_27_29 ( .A(u5_mult_82_ab_27__29_), .B(
        u5_mult_82_CARRYB_26__29_), .CI(u5_mult_82_SUMB_26__30_), .CO(
        u5_mult_82_CARRYB_27__29_), .S(u5_mult_82_SUMB_27__29_) );
  FA_X1 u5_mult_82_S2_27_28 ( .A(u5_mult_82_ab_27__28_), .B(
        u5_mult_82_CARRYB_26__28_), .CI(u5_mult_82_SUMB_26__29_), .CO(
        u5_mult_82_CARRYB_27__28_), .S(u5_mult_82_SUMB_27__28_) );
  FA_X1 u5_mult_82_S2_27_27 ( .A(u5_mult_82_ab_27__27_), .B(
        u5_mult_82_CARRYB_26__27_), .CI(u5_mult_82_SUMB_26__28_), .CO(
        u5_mult_82_CARRYB_27__27_), .S(u5_mult_82_SUMB_27__27_) );
  FA_X1 u5_mult_82_S2_27_26 ( .A(u5_mult_82_ab_27__26_), .B(
        u5_mult_82_CARRYB_26__26_), .CI(u5_mult_82_SUMB_26__27_), .CO(
        u5_mult_82_CARRYB_27__26_), .S(u5_mult_82_SUMB_27__26_) );
  FA_X1 u5_mult_82_S2_27_25 ( .A(u5_mult_82_ab_27__25_), .B(
        u5_mult_82_CARRYB_26__25_), .CI(u5_mult_82_SUMB_26__26_), .CO(
        u5_mult_82_CARRYB_27__25_), .S(u5_mult_82_SUMB_27__25_) );
  FA_X1 u5_mult_82_S2_27_24 ( .A(u5_mult_82_ab_27__24_), .B(
        u5_mult_82_CARRYB_26__24_), .CI(u5_mult_82_SUMB_26__25_), .CO(
        u5_mult_82_CARRYB_27__24_), .S(u5_mult_82_SUMB_27__24_) );
  FA_X1 u5_mult_82_S2_27_23 ( .A(u5_mult_82_ab_27__23_), .B(
        u5_mult_82_CARRYB_26__23_), .CI(u5_mult_82_SUMB_26__24_), .CO(
        u5_mult_82_CARRYB_27__23_), .S(u5_mult_82_SUMB_27__23_) );
  FA_X1 u5_mult_82_S2_27_22 ( .A(u5_mult_82_ab_27__22_), .B(
        u5_mult_82_CARRYB_26__22_), .CI(u5_mult_82_SUMB_26__23_), .CO(
        u5_mult_82_CARRYB_27__22_), .S(u5_mult_82_SUMB_27__22_) );
  FA_X1 u5_mult_82_S2_27_21 ( .A(u5_mult_82_ab_27__21_), .B(
        u5_mult_82_CARRYB_26__21_), .CI(u5_mult_82_SUMB_26__22_), .CO(
        u5_mult_82_CARRYB_27__21_), .S(u5_mult_82_SUMB_27__21_) );
  FA_X1 u5_mult_82_S2_27_20 ( .A(u5_mult_82_ab_27__20_), .B(
        u5_mult_82_CARRYB_26__20_), .CI(u5_mult_82_SUMB_26__21_), .CO(
        u5_mult_82_CARRYB_27__20_), .S(u5_mult_82_SUMB_27__20_) );
  FA_X1 u5_mult_82_S2_27_19 ( .A(u5_mult_82_ab_27__19_), .B(
        u5_mult_82_CARRYB_26__19_), .CI(u5_mult_82_SUMB_26__20_), .CO(
        u5_mult_82_CARRYB_27__19_), .S(u5_mult_82_SUMB_27__19_) );
  FA_X1 u5_mult_82_S2_27_18 ( .A(u5_mult_82_ab_27__18_), .B(
        u5_mult_82_CARRYB_26__18_), .CI(u5_mult_82_SUMB_26__19_), .CO(
        u5_mult_82_CARRYB_27__18_), .S(u5_mult_82_SUMB_27__18_) );
  FA_X1 u5_mult_82_S2_27_17 ( .A(u5_mult_82_ab_27__17_), .B(
        u5_mult_82_CARRYB_26__17_), .CI(u5_mult_82_SUMB_26__18_), .CO(
        u5_mult_82_CARRYB_27__17_), .S(u5_mult_82_SUMB_27__17_) );
  FA_X1 u5_mult_82_S2_27_16 ( .A(u5_mult_82_ab_27__16_), .B(
        u5_mult_82_CARRYB_26__16_), .CI(u5_mult_82_SUMB_26__17_), .CO(
        u5_mult_82_CARRYB_27__16_), .S(u5_mult_82_SUMB_27__16_) );
  FA_X1 u5_mult_82_S2_27_15 ( .A(u5_mult_82_ab_27__15_), .B(
        u5_mult_82_CARRYB_26__15_), .CI(u5_mult_82_SUMB_26__16_), .CO(
        u5_mult_82_CARRYB_27__15_), .S(u5_mult_82_SUMB_27__15_) );
  FA_X1 u5_mult_82_S2_27_14 ( .A(u5_mult_82_ab_27__14_), .B(
        u5_mult_82_CARRYB_26__14_), .CI(u5_mult_82_SUMB_26__15_), .CO(
        u5_mult_82_CARRYB_27__14_), .S(u5_mult_82_SUMB_27__14_) );
  FA_X1 u5_mult_82_S2_27_13 ( .A(u5_mult_82_ab_27__13_), .B(
        u5_mult_82_CARRYB_26__13_), .CI(u5_mult_82_SUMB_26__14_), .CO(
        u5_mult_82_CARRYB_27__13_), .S(u5_mult_82_SUMB_27__13_) );
  FA_X1 u5_mult_82_S2_27_12 ( .A(u5_mult_82_ab_27__12_), .B(
        u5_mult_82_CARRYB_26__12_), .CI(u5_mult_82_SUMB_26__13_), .CO(
        u5_mult_82_CARRYB_27__12_), .S(u5_mult_82_SUMB_27__12_) );
  FA_X1 u5_mult_82_S2_27_11 ( .A(u5_mult_82_ab_27__11_), .B(
        u5_mult_82_CARRYB_26__11_), .CI(u5_mult_82_SUMB_26__12_), .CO(
        u5_mult_82_CARRYB_27__11_), .S(u5_mult_82_SUMB_27__11_) );
  FA_X1 u5_mult_82_S2_27_10 ( .A(u5_mult_82_ab_27__10_), .B(
        u5_mult_82_CARRYB_26__10_), .CI(u5_mult_82_SUMB_26__11_), .CO(
        u5_mult_82_CARRYB_27__10_), .S(u5_mult_82_SUMB_27__10_) );
  FA_X1 u5_mult_82_S2_27_9 ( .A(u5_mult_82_ab_27__9_), .B(
        u5_mult_82_CARRYB_26__9_), .CI(u5_mult_82_SUMB_26__10_), .CO(
        u5_mult_82_CARRYB_27__9_), .S(u5_mult_82_SUMB_27__9_) );
  FA_X1 u5_mult_82_S2_27_8 ( .A(u5_mult_82_ab_27__8_), .B(
        u5_mult_82_CARRYB_26__8_), .CI(u5_mult_82_SUMB_26__9_), .CO(
        u5_mult_82_CARRYB_27__8_), .S(u5_mult_82_SUMB_27__8_) );
  FA_X1 u5_mult_82_S2_27_7 ( .A(u5_mult_82_ab_27__7_), .B(
        u5_mult_82_CARRYB_26__7_), .CI(u5_mult_82_SUMB_26__8_), .CO(
        u5_mult_82_CARRYB_27__7_), .S(u5_mult_82_SUMB_27__7_) );
  FA_X1 u5_mult_82_S2_27_6 ( .A(u5_mult_82_ab_27__6_), .B(
        u5_mult_82_CARRYB_26__6_), .CI(u5_mult_82_SUMB_26__7_), .CO(
        u5_mult_82_CARRYB_27__6_), .S(u5_mult_82_SUMB_27__6_) );
  FA_X1 u5_mult_82_S2_27_5 ( .A(u5_mult_82_ab_27__5_), .B(
        u5_mult_82_CARRYB_26__5_), .CI(u5_mult_82_SUMB_26__6_), .CO(
        u5_mult_82_CARRYB_27__5_), .S(u5_mult_82_SUMB_27__5_) );
  FA_X1 u5_mult_82_S2_27_4 ( .A(u5_mult_82_ab_27__4_), .B(
        u5_mult_82_CARRYB_26__4_), .CI(u5_mult_82_SUMB_26__5_), .CO(
        u5_mult_82_CARRYB_27__4_), .S(u5_mult_82_SUMB_27__4_) );
  FA_X1 u5_mult_82_S2_27_3 ( .A(u5_mult_82_ab_27__3_), .B(
        u5_mult_82_CARRYB_26__3_), .CI(u5_mult_82_SUMB_26__4_), .CO(
        u5_mult_82_CARRYB_27__3_), .S(u5_mult_82_SUMB_27__3_) );
  FA_X1 u5_mult_82_S2_27_2 ( .A(u5_mult_82_ab_27__2_), .B(
        u5_mult_82_CARRYB_26__2_), .CI(u5_mult_82_SUMB_26__3_), .CO(
        u5_mult_82_CARRYB_27__2_), .S(u5_mult_82_SUMB_27__2_) );
  FA_X1 u5_mult_82_S2_27_1 ( .A(u5_mult_82_ab_27__1_), .B(
        u5_mult_82_CARRYB_26__1_), .CI(u5_mult_82_SUMB_26__2_), .CO(
        u5_mult_82_CARRYB_27__1_), .S(u5_mult_82_SUMB_27__1_) );
  FA_X1 u5_mult_82_S1_27_0 ( .A(u5_mult_82_ab_27__0_), .B(
        u5_mult_82_CARRYB_26__0_), .CI(u5_mult_82_SUMB_26__1_), .CO(
        u5_mult_82_CARRYB_27__0_), .S(u5_N27) );
  FA_X1 u5_mult_82_S3_28_51 ( .A(u5_mult_82_ab_28__51_), .B(
        u5_mult_82_CARRYB_27__51_), .CI(u5_mult_82_ab_27__52_), .CO(
        u5_mult_82_CARRYB_28__51_), .S(u5_mult_82_SUMB_28__51_) );
  FA_X1 u5_mult_82_S2_28_50 ( .A(u5_mult_82_ab_28__50_), .B(
        u5_mult_82_CARRYB_27__50_), .CI(u5_mult_82_SUMB_27__51_), .CO(
        u5_mult_82_CARRYB_28__50_), .S(u5_mult_82_SUMB_28__50_) );
  FA_X1 u5_mult_82_S2_28_49 ( .A(u5_mult_82_ab_28__49_), .B(
        u5_mult_82_CARRYB_27__49_), .CI(u5_mult_82_SUMB_27__50_), .CO(
        u5_mult_82_CARRYB_28__49_), .S(u5_mult_82_SUMB_28__49_) );
  FA_X1 u5_mult_82_S2_28_48 ( .A(u5_mult_82_ab_28__48_), .B(
        u5_mult_82_CARRYB_27__48_), .CI(u5_mult_82_SUMB_27__49_), .CO(
        u5_mult_82_CARRYB_28__48_), .S(u5_mult_82_SUMB_28__48_) );
  FA_X1 u5_mult_82_S2_28_47 ( .A(u5_mult_82_ab_28__47_), .B(
        u5_mult_82_CARRYB_27__47_), .CI(u5_mult_82_SUMB_27__48_), .CO(
        u5_mult_82_CARRYB_28__47_), .S(u5_mult_82_SUMB_28__47_) );
  FA_X1 u5_mult_82_S2_28_46 ( .A(u5_mult_82_ab_28__46_), .B(
        u5_mult_82_CARRYB_27__46_), .CI(u5_mult_82_SUMB_27__47_), .CO(
        u5_mult_82_CARRYB_28__46_), .S(u5_mult_82_SUMB_28__46_) );
  FA_X1 u5_mult_82_S2_28_45 ( .A(u5_mult_82_ab_28__45_), .B(
        u5_mult_82_CARRYB_27__45_), .CI(u5_mult_82_SUMB_27__46_), .CO(
        u5_mult_82_CARRYB_28__45_), .S(u5_mult_82_SUMB_28__45_) );
  FA_X1 u5_mult_82_S2_28_44 ( .A(u5_mult_82_ab_28__44_), .B(
        u5_mult_82_CARRYB_27__44_), .CI(u5_mult_82_SUMB_27__45_), .CO(
        u5_mult_82_CARRYB_28__44_), .S(u5_mult_82_SUMB_28__44_) );
  FA_X1 u5_mult_82_S2_28_43 ( .A(u5_mult_82_ab_28__43_), .B(
        u5_mult_82_CARRYB_27__43_), .CI(u5_mult_82_SUMB_27__44_), .CO(
        u5_mult_82_CARRYB_28__43_), .S(u5_mult_82_SUMB_28__43_) );
  FA_X1 u5_mult_82_S2_28_42 ( .A(u5_mult_82_ab_28__42_), .B(
        u5_mult_82_CARRYB_27__42_), .CI(u5_mult_82_SUMB_27__43_), .CO(
        u5_mult_82_CARRYB_28__42_), .S(u5_mult_82_SUMB_28__42_) );
  FA_X1 u5_mult_82_S2_28_41 ( .A(u5_mult_82_ab_28__41_), .B(
        u5_mult_82_CARRYB_27__41_), .CI(u5_mult_82_SUMB_27__42_), .CO(
        u5_mult_82_CARRYB_28__41_), .S(u5_mult_82_SUMB_28__41_) );
  FA_X1 u5_mult_82_S2_28_40 ( .A(u5_mult_82_ab_28__40_), .B(
        u5_mult_82_CARRYB_27__40_), .CI(u5_mult_82_SUMB_27__41_), .CO(
        u5_mult_82_CARRYB_28__40_), .S(u5_mult_82_SUMB_28__40_) );
  FA_X1 u5_mult_82_S2_28_39 ( .A(u5_mult_82_ab_28__39_), .B(
        u5_mult_82_CARRYB_27__39_), .CI(u5_mult_82_SUMB_27__40_), .CO(
        u5_mult_82_CARRYB_28__39_), .S(u5_mult_82_SUMB_28__39_) );
  FA_X1 u5_mult_82_S2_28_38 ( .A(u5_mult_82_ab_28__38_), .B(
        u5_mult_82_CARRYB_27__38_), .CI(u5_mult_82_SUMB_27__39_), .CO(
        u5_mult_82_CARRYB_28__38_), .S(u5_mult_82_SUMB_28__38_) );
  FA_X1 u5_mult_82_S2_28_37 ( .A(u5_mult_82_ab_28__37_), .B(
        u5_mult_82_CARRYB_27__37_), .CI(u5_mult_82_SUMB_27__38_), .CO(
        u5_mult_82_CARRYB_28__37_), .S(u5_mult_82_SUMB_28__37_) );
  FA_X1 u5_mult_82_S2_28_36 ( .A(u5_mult_82_ab_28__36_), .B(
        u5_mult_82_CARRYB_27__36_), .CI(u5_mult_82_SUMB_27__37_), .CO(
        u5_mult_82_CARRYB_28__36_), .S(u5_mult_82_SUMB_28__36_) );
  FA_X1 u5_mult_82_S2_28_35 ( .A(u5_mult_82_ab_28__35_), .B(
        u5_mult_82_CARRYB_27__35_), .CI(u5_mult_82_SUMB_27__36_), .CO(
        u5_mult_82_CARRYB_28__35_), .S(u5_mult_82_SUMB_28__35_) );
  FA_X1 u5_mult_82_S2_28_34 ( .A(u5_mult_82_ab_28__34_), .B(
        u5_mult_82_CARRYB_27__34_), .CI(u5_mult_82_SUMB_27__35_), .CO(
        u5_mult_82_CARRYB_28__34_), .S(u5_mult_82_SUMB_28__34_) );
  FA_X1 u5_mult_82_S2_28_33 ( .A(u5_mult_82_ab_28__33_), .B(
        u5_mult_82_CARRYB_27__33_), .CI(u5_mult_82_SUMB_27__34_), .CO(
        u5_mult_82_CARRYB_28__33_), .S(u5_mult_82_SUMB_28__33_) );
  FA_X1 u5_mult_82_S2_28_32 ( .A(u5_mult_82_ab_28__32_), .B(
        u5_mult_82_CARRYB_27__32_), .CI(u5_mult_82_SUMB_27__33_), .CO(
        u5_mult_82_CARRYB_28__32_), .S(u5_mult_82_SUMB_28__32_) );
  FA_X1 u5_mult_82_S2_28_31 ( .A(u5_mult_82_ab_28__31_), .B(
        u5_mult_82_CARRYB_27__31_), .CI(u5_mult_82_SUMB_27__32_), .CO(
        u5_mult_82_CARRYB_28__31_), .S(u5_mult_82_SUMB_28__31_) );
  FA_X1 u5_mult_82_S2_28_30 ( .A(u5_mult_82_ab_28__30_), .B(
        u5_mult_82_CARRYB_27__30_), .CI(u5_mult_82_SUMB_27__31_), .CO(
        u5_mult_82_CARRYB_28__30_), .S(u5_mult_82_SUMB_28__30_) );
  FA_X1 u5_mult_82_S2_28_29 ( .A(u5_mult_82_ab_28__29_), .B(
        u5_mult_82_CARRYB_27__29_), .CI(u5_mult_82_SUMB_27__30_), .CO(
        u5_mult_82_CARRYB_28__29_), .S(u5_mult_82_SUMB_28__29_) );
  FA_X1 u5_mult_82_S2_28_28 ( .A(u5_mult_82_ab_28__28_), .B(
        u5_mult_82_CARRYB_27__28_), .CI(u5_mult_82_SUMB_27__29_), .CO(
        u5_mult_82_CARRYB_28__28_), .S(u5_mult_82_SUMB_28__28_) );
  FA_X1 u5_mult_82_S2_28_27 ( .A(u5_mult_82_ab_28__27_), .B(
        u5_mult_82_CARRYB_27__27_), .CI(u5_mult_82_SUMB_27__28_), .CO(
        u5_mult_82_CARRYB_28__27_), .S(u5_mult_82_SUMB_28__27_) );
  FA_X1 u5_mult_82_S2_28_26 ( .A(u5_mult_82_ab_28__26_), .B(
        u5_mult_82_CARRYB_27__26_), .CI(u5_mult_82_SUMB_27__27_), .CO(
        u5_mult_82_CARRYB_28__26_), .S(u5_mult_82_SUMB_28__26_) );
  FA_X1 u5_mult_82_S2_28_25 ( .A(u5_mult_82_ab_28__25_), .B(
        u5_mult_82_CARRYB_27__25_), .CI(u5_mult_82_SUMB_27__26_), .CO(
        u5_mult_82_CARRYB_28__25_), .S(u5_mult_82_SUMB_28__25_) );
  FA_X1 u5_mult_82_S2_28_24 ( .A(u5_mult_82_ab_28__24_), .B(
        u5_mult_82_CARRYB_27__24_), .CI(u5_mult_82_SUMB_27__25_), .CO(
        u5_mult_82_CARRYB_28__24_), .S(u5_mult_82_SUMB_28__24_) );
  FA_X1 u5_mult_82_S2_28_23 ( .A(u5_mult_82_ab_28__23_), .B(
        u5_mult_82_CARRYB_27__23_), .CI(u5_mult_82_SUMB_27__24_), .CO(
        u5_mult_82_CARRYB_28__23_), .S(u5_mult_82_SUMB_28__23_) );
  FA_X1 u5_mult_82_S2_28_22 ( .A(u5_mult_82_ab_28__22_), .B(
        u5_mult_82_CARRYB_27__22_), .CI(u5_mult_82_SUMB_27__23_), .CO(
        u5_mult_82_CARRYB_28__22_), .S(u5_mult_82_SUMB_28__22_) );
  FA_X1 u5_mult_82_S2_28_21 ( .A(u5_mult_82_ab_28__21_), .B(
        u5_mult_82_CARRYB_27__21_), .CI(u5_mult_82_SUMB_27__22_), .CO(
        u5_mult_82_CARRYB_28__21_), .S(u5_mult_82_SUMB_28__21_) );
  FA_X1 u5_mult_82_S2_28_20 ( .A(u5_mult_82_ab_28__20_), .B(
        u5_mult_82_CARRYB_27__20_), .CI(u5_mult_82_SUMB_27__21_), .CO(
        u5_mult_82_CARRYB_28__20_), .S(u5_mult_82_SUMB_28__20_) );
  FA_X1 u5_mult_82_S2_28_19 ( .A(u5_mult_82_ab_28__19_), .B(
        u5_mult_82_CARRYB_27__19_), .CI(u5_mult_82_SUMB_27__20_), .CO(
        u5_mult_82_CARRYB_28__19_), .S(u5_mult_82_SUMB_28__19_) );
  FA_X1 u5_mult_82_S2_28_18 ( .A(u5_mult_82_ab_28__18_), .B(
        u5_mult_82_CARRYB_27__18_), .CI(u5_mult_82_SUMB_27__19_), .CO(
        u5_mult_82_CARRYB_28__18_), .S(u5_mult_82_SUMB_28__18_) );
  FA_X1 u5_mult_82_S2_28_17 ( .A(u5_mult_82_ab_28__17_), .B(
        u5_mult_82_CARRYB_27__17_), .CI(u5_mult_82_SUMB_27__18_), .CO(
        u5_mult_82_CARRYB_28__17_), .S(u5_mult_82_SUMB_28__17_) );
  FA_X1 u5_mult_82_S2_28_16 ( .A(u5_mult_82_ab_28__16_), .B(
        u5_mult_82_CARRYB_27__16_), .CI(u5_mult_82_SUMB_27__17_), .CO(
        u5_mult_82_CARRYB_28__16_), .S(u5_mult_82_SUMB_28__16_) );
  FA_X1 u5_mult_82_S2_28_15 ( .A(u5_mult_82_ab_28__15_), .B(
        u5_mult_82_CARRYB_27__15_), .CI(u5_mult_82_SUMB_27__16_), .CO(
        u5_mult_82_CARRYB_28__15_), .S(u5_mult_82_SUMB_28__15_) );
  FA_X1 u5_mult_82_S2_28_14 ( .A(u5_mult_82_ab_28__14_), .B(
        u5_mult_82_CARRYB_27__14_), .CI(u5_mult_82_SUMB_27__15_), .CO(
        u5_mult_82_CARRYB_28__14_), .S(u5_mult_82_SUMB_28__14_) );
  FA_X1 u5_mult_82_S2_28_13 ( .A(u5_mult_82_ab_28__13_), .B(
        u5_mult_82_CARRYB_27__13_), .CI(u5_mult_82_SUMB_27__14_), .CO(
        u5_mult_82_CARRYB_28__13_), .S(u5_mult_82_SUMB_28__13_) );
  FA_X1 u5_mult_82_S2_28_12 ( .A(u5_mult_82_ab_28__12_), .B(
        u5_mult_82_CARRYB_27__12_), .CI(u5_mult_82_SUMB_27__13_), .CO(
        u5_mult_82_CARRYB_28__12_), .S(u5_mult_82_SUMB_28__12_) );
  FA_X1 u5_mult_82_S2_28_11 ( .A(u5_mult_82_ab_28__11_), .B(
        u5_mult_82_CARRYB_27__11_), .CI(u5_mult_82_SUMB_27__12_), .CO(
        u5_mult_82_CARRYB_28__11_), .S(u5_mult_82_SUMB_28__11_) );
  FA_X1 u5_mult_82_S2_28_10 ( .A(u5_mult_82_ab_28__10_), .B(
        u5_mult_82_CARRYB_27__10_), .CI(u5_mult_82_SUMB_27__11_), .CO(
        u5_mult_82_CARRYB_28__10_), .S(u5_mult_82_SUMB_28__10_) );
  FA_X1 u5_mult_82_S2_28_9 ( .A(u5_mult_82_ab_28__9_), .B(
        u5_mult_82_CARRYB_27__9_), .CI(u5_mult_82_SUMB_27__10_), .CO(
        u5_mult_82_CARRYB_28__9_), .S(u5_mult_82_SUMB_28__9_) );
  FA_X1 u5_mult_82_S2_28_8 ( .A(u5_mult_82_ab_28__8_), .B(
        u5_mult_82_CARRYB_27__8_), .CI(u5_mult_82_SUMB_27__9_), .CO(
        u5_mult_82_CARRYB_28__8_), .S(u5_mult_82_SUMB_28__8_) );
  FA_X1 u5_mult_82_S2_28_7 ( .A(u5_mult_82_ab_28__7_), .B(
        u5_mult_82_CARRYB_27__7_), .CI(u5_mult_82_SUMB_27__8_), .CO(
        u5_mult_82_CARRYB_28__7_), .S(u5_mult_82_SUMB_28__7_) );
  FA_X1 u5_mult_82_S2_28_6 ( .A(u5_mult_82_ab_28__6_), .B(
        u5_mult_82_CARRYB_27__6_), .CI(u5_mult_82_SUMB_27__7_), .CO(
        u5_mult_82_CARRYB_28__6_), .S(u5_mult_82_SUMB_28__6_) );
  FA_X1 u5_mult_82_S2_28_5 ( .A(u5_mult_82_ab_28__5_), .B(
        u5_mult_82_CARRYB_27__5_), .CI(u5_mult_82_SUMB_27__6_), .CO(
        u5_mult_82_CARRYB_28__5_), .S(u5_mult_82_SUMB_28__5_) );
  FA_X1 u5_mult_82_S2_28_4 ( .A(u5_mult_82_ab_28__4_), .B(
        u5_mult_82_CARRYB_27__4_), .CI(u5_mult_82_SUMB_27__5_), .CO(
        u5_mult_82_CARRYB_28__4_), .S(u5_mult_82_SUMB_28__4_) );
  FA_X1 u5_mult_82_S2_28_3 ( .A(u5_mult_82_ab_28__3_), .B(
        u5_mult_82_CARRYB_27__3_), .CI(u5_mult_82_SUMB_27__4_), .CO(
        u5_mult_82_CARRYB_28__3_), .S(u5_mult_82_SUMB_28__3_) );
  FA_X1 u5_mult_82_S2_28_2 ( .A(u5_mult_82_ab_28__2_), .B(
        u5_mult_82_CARRYB_27__2_), .CI(u5_mult_82_SUMB_27__3_), .CO(
        u5_mult_82_CARRYB_28__2_), .S(u5_mult_82_SUMB_28__2_) );
  FA_X1 u5_mult_82_S2_28_1 ( .A(u5_mult_82_ab_28__1_), .B(
        u5_mult_82_CARRYB_27__1_), .CI(u5_mult_82_SUMB_27__2_), .CO(
        u5_mult_82_CARRYB_28__1_), .S(u5_mult_82_SUMB_28__1_) );
  FA_X1 u5_mult_82_S1_28_0 ( .A(u5_mult_82_ab_28__0_), .B(
        u5_mult_82_CARRYB_27__0_), .CI(u5_mult_82_SUMB_27__1_), .CO(
        u5_mult_82_CARRYB_28__0_), .S(u5_N28) );
  FA_X1 u5_mult_82_S3_29_51 ( .A(u5_mult_82_ab_29__51_), .B(
        u5_mult_82_CARRYB_28__51_), .CI(u5_mult_82_ab_28__52_), .CO(
        u5_mult_82_CARRYB_29__51_), .S(u5_mult_82_SUMB_29__51_) );
  FA_X1 u5_mult_82_S2_29_50 ( .A(u5_mult_82_ab_29__50_), .B(
        u5_mult_82_CARRYB_28__50_), .CI(u5_mult_82_SUMB_28__51_), .CO(
        u5_mult_82_CARRYB_29__50_), .S(u5_mult_82_SUMB_29__50_) );
  FA_X1 u5_mult_82_S2_29_49 ( .A(u5_mult_82_ab_29__49_), .B(
        u5_mult_82_CARRYB_28__49_), .CI(u5_mult_82_SUMB_28__50_), .CO(
        u5_mult_82_CARRYB_29__49_), .S(u5_mult_82_SUMB_29__49_) );
  FA_X1 u5_mult_82_S2_29_48 ( .A(u5_mult_82_ab_29__48_), .B(
        u5_mult_82_CARRYB_28__48_), .CI(u5_mult_82_SUMB_28__49_), .CO(
        u5_mult_82_CARRYB_29__48_), .S(u5_mult_82_SUMB_29__48_) );
  FA_X1 u5_mult_82_S2_29_47 ( .A(u5_mult_82_ab_29__47_), .B(
        u5_mult_82_CARRYB_28__47_), .CI(u5_mult_82_SUMB_28__48_), .CO(
        u5_mult_82_CARRYB_29__47_), .S(u5_mult_82_SUMB_29__47_) );
  FA_X1 u5_mult_82_S2_29_46 ( .A(u5_mult_82_ab_29__46_), .B(
        u5_mult_82_CARRYB_28__46_), .CI(u5_mult_82_SUMB_28__47_), .CO(
        u5_mult_82_CARRYB_29__46_), .S(u5_mult_82_SUMB_29__46_) );
  FA_X1 u5_mult_82_S2_29_45 ( .A(u5_mult_82_ab_29__45_), .B(
        u5_mult_82_CARRYB_28__45_), .CI(u5_mult_82_SUMB_28__46_), .CO(
        u5_mult_82_CARRYB_29__45_), .S(u5_mult_82_SUMB_29__45_) );
  FA_X1 u5_mult_82_S2_29_44 ( .A(u5_mult_82_ab_29__44_), .B(
        u5_mult_82_CARRYB_28__44_), .CI(u5_mult_82_SUMB_28__45_), .CO(
        u5_mult_82_CARRYB_29__44_), .S(u5_mult_82_SUMB_29__44_) );
  FA_X1 u5_mult_82_S2_29_43 ( .A(u5_mult_82_ab_29__43_), .B(
        u5_mult_82_CARRYB_28__43_), .CI(u5_mult_82_SUMB_28__44_), .CO(
        u5_mult_82_CARRYB_29__43_), .S(u5_mult_82_SUMB_29__43_) );
  FA_X1 u5_mult_82_S2_29_42 ( .A(u5_mult_82_ab_29__42_), .B(
        u5_mult_82_CARRYB_28__42_), .CI(u5_mult_82_SUMB_28__43_), .CO(
        u5_mult_82_CARRYB_29__42_), .S(u5_mult_82_SUMB_29__42_) );
  FA_X1 u5_mult_82_S2_29_41 ( .A(u5_mult_82_ab_29__41_), .B(
        u5_mult_82_CARRYB_28__41_), .CI(u5_mult_82_SUMB_28__42_), .CO(
        u5_mult_82_CARRYB_29__41_), .S(u5_mult_82_SUMB_29__41_) );
  FA_X1 u5_mult_82_S2_29_40 ( .A(u5_mult_82_ab_29__40_), .B(
        u5_mult_82_CARRYB_28__40_), .CI(u5_mult_82_SUMB_28__41_), .CO(
        u5_mult_82_CARRYB_29__40_), .S(u5_mult_82_SUMB_29__40_) );
  FA_X1 u5_mult_82_S2_29_39 ( .A(u5_mult_82_ab_29__39_), .B(
        u5_mult_82_CARRYB_28__39_), .CI(u5_mult_82_SUMB_28__40_), .CO(
        u5_mult_82_CARRYB_29__39_), .S(u5_mult_82_SUMB_29__39_) );
  FA_X1 u5_mult_82_S2_29_38 ( .A(u5_mult_82_ab_29__38_), .B(
        u5_mult_82_CARRYB_28__38_), .CI(u5_mult_82_SUMB_28__39_), .CO(
        u5_mult_82_CARRYB_29__38_), .S(u5_mult_82_SUMB_29__38_) );
  FA_X1 u5_mult_82_S2_29_37 ( .A(u5_mult_82_ab_29__37_), .B(
        u5_mult_82_CARRYB_28__37_), .CI(u5_mult_82_SUMB_28__38_), .CO(
        u5_mult_82_CARRYB_29__37_), .S(u5_mult_82_SUMB_29__37_) );
  FA_X1 u5_mult_82_S2_29_36 ( .A(u5_mult_82_ab_29__36_), .B(
        u5_mult_82_CARRYB_28__36_), .CI(u5_mult_82_SUMB_28__37_), .CO(
        u5_mult_82_CARRYB_29__36_), .S(u5_mult_82_SUMB_29__36_) );
  FA_X1 u5_mult_82_S2_29_35 ( .A(u5_mult_82_ab_29__35_), .B(
        u5_mult_82_CARRYB_28__35_), .CI(u5_mult_82_SUMB_28__36_), .CO(
        u5_mult_82_CARRYB_29__35_), .S(u5_mult_82_SUMB_29__35_) );
  FA_X1 u5_mult_82_S2_29_34 ( .A(u5_mult_82_ab_29__34_), .B(
        u5_mult_82_CARRYB_28__34_), .CI(u5_mult_82_SUMB_28__35_), .CO(
        u5_mult_82_CARRYB_29__34_), .S(u5_mult_82_SUMB_29__34_) );
  FA_X1 u5_mult_82_S2_29_33 ( .A(u5_mult_82_ab_29__33_), .B(
        u5_mult_82_CARRYB_28__33_), .CI(u5_mult_82_SUMB_28__34_), .CO(
        u5_mult_82_CARRYB_29__33_), .S(u5_mult_82_SUMB_29__33_) );
  FA_X1 u5_mult_82_S2_29_32 ( .A(u5_mult_82_ab_29__32_), .B(
        u5_mult_82_CARRYB_28__32_), .CI(u5_mult_82_SUMB_28__33_), .CO(
        u5_mult_82_CARRYB_29__32_), .S(u5_mult_82_SUMB_29__32_) );
  FA_X1 u5_mult_82_S2_29_31 ( .A(u5_mult_82_ab_29__31_), .B(
        u5_mult_82_CARRYB_28__31_), .CI(u5_mult_82_SUMB_28__32_), .CO(
        u5_mult_82_CARRYB_29__31_), .S(u5_mult_82_SUMB_29__31_) );
  FA_X1 u5_mult_82_S2_29_30 ( .A(u5_mult_82_ab_29__30_), .B(
        u5_mult_82_CARRYB_28__30_), .CI(u5_mult_82_SUMB_28__31_), .CO(
        u5_mult_82_CARRYB_29__30_), .S(u5_mult_82_SUMB_29__30_) );
  FA_X1 u5_mult_82_S2_29_29 ( .A(u5_mult_82_ab_29__29_), .B(
        u5_mult_82_CARRYB_28__29_), .CI(u5_mult_82_SUMB_28__30_), .CO(
        u5_mult_82_CARRYB_29__29_), .S(u5_mult_82_SUMB_29__29_) );
  FA_X1 u5_mult_82_S2_29_28 ( .A(u5_mult_82_ab_29__28_), .B(
        u5_mult_82_CARRYB_28__28_), .CI(u5_mult_82_SUMB_28__29_), .CO(
        u5_mult_82_CARRYB_29__28_), .S(u5_mult_82_SUMB_29__28_) );
  FA_X1 u5_mult_82_S2_29_27 ( .A(u5_mult_82_ab_29__27_), .B(
        u5_mult_82_CARRYB_28__27_), .CI(u5_mult_82_SUMB_28__28_), .CO(
        u5_mult_82_CARRYB_29__27_), .S(u5_mult_82_SUMB_29__27_) );
  FA_X1 u5_mult_82_S2_29_26 ( .A(u5_mult_82_ab_29__26_), .B(
        u5_mult_82_CARRYB_28__26_), .CI(u5_mult_82_SUMB_28__27_), .CO(
        u5_mult_82_CARRYB_29__26_), .S(u5_mult_82_SUMB_29__26_) );
  FA_X1 u5_mult_82_S2_29_25 ( .A(u5_mult_82_ab_29__25_), .B(
        u5_mult_82_CARRYB_28__25_), .CI(u5_mult_82_SUMB_28__26_), .CO(
        u5_mult_82_CARRYB_29__25_), .S(u5_mult_82_SUMB_29__25_) );
  FA_X1 u5_mult_82_S2_29_24 ( .A(u5_mult_82_ab_29__24_), .B(
        u5_mult_82_CARRYB_28__24_), .CI(u5_mult_82_SUMB_28__25_), .CO(
        u5_mult_82_CARRYB_29__24_), .S(u5_mult_82_SUMB_29__24_) );
  FA_X1 u5_mult_82_S2_29_23 ( .A(u5_mult_82_ab_29__23_), .B(
        u5_mult_82_CARRYB_28__23_), .CI(u5_mult_82_SUMB_28__24_), .CO(
        u5_mult_82_CARRYB_29__23_), .S(u5_mult_82_SUMB_29__23_) );
  FA_X1 u5_mult_82_S2_29_22 ( .A(u5_mult_82_ab_29__22_), .B(
        u5_mult_82_CARRYB_28__22_), .CI(u5_mult_82_SUMB_28__23_), .CO(
        u5_mult_82_CARRYB_29__22_), .S(u5_mult_82_SUMB_29__22_) );
  FA_X1 u5_mult_82_S2_29_21 ( .A(u5_mult_82_ab_29__21_), .B(
        u5_mult_82_CARRYB_28__21_), .CI(u5_mult_82_SUMB_28__22_), .CO(
        u5_mult_82_CARRYB_29__21_), .S(u5_mult_82_SUMB_29__21_) );
  FA_X1 u5_mult_82_S2_29_20 ( .A(u5_mult_82_ab_29__20_), .B(
        u5_mult_82_CARRYB_28__20_), .CI(u5_mult_82_SUMB_28__21_), .CO(
        u5_mult_82_CARRYB_29__20_), .S(u5_mult_82_SUMB_29__20_) );
  FA_X1 u5_mult_82_S2_29_19 ( .A(u5_mult_82_ab_29__19_), .B(
        u5_mult_82_CARRYB_28__19_), .CI(u5_mult_82_SUMB_28__20_), .CO(
        u5_mult_82_CARRYB_29__19_), .S(u5_mult_82_SUMB_29__19_) );
  FA_X1 u5_mult_82_S2_29_18 ( .A(u5_mult_82_ab_29__18_), .B(
        u5_mult_82_CARRYB_28__18_), .CI(u5_mult_82_SUMB_28__19_), .CO(
        u5_mult_82_CARRYB_29__18_), .S(u5_mult_82_SUMB_29__18_) );
  FA_X1 u5_mult_82_S2_29_17 ( .A(u5_mult_82_ab_29__17_), .B(
        u5_mult_82_CARRYB_28__17_), .CI(u5_mult_82_SUMB_28__18_), .CO(
        u5_mult_82_CARRYB_29__17_), .S(u5_mult_82_SUMB_29__17_) );
  FA_X1 u5_mult_82_S2_29_16 ( .A(u5_mult_82_ab_29__16_), .B(
        u5_mult_82_CARRYB_28__16_), .CI(u5_mult_82_SUMB_28__17_), .CO(
        u5_mult_82_CARRYB_29__16_), .S(u5_mult_82_SUMB_29__16_) );
  FA_X1 u5_mult_82_S2_29_15 ( .A(u5_mult_82_ab_29__15_), .B(
        u5_mult_82_CARRYB_28__15_), .CI(u5_mult_82_SUMB_28__16_), .CO(
        u5_mult_82_CARRYB_29__15_), .S(u5_mult_82_SUMB_29__15_) );
  FA_X1 u5_mult_82_S2_29_14 ( .A(u5_mult_82_ab_29__14_), .B(
        u5_mult_82_CARRYB_28__14_), .CI(u5_mult_82_SUMB_28__15_), .CO(
        u5_mult_82_CARRYB_29__14_), .S(u5_mult_82_SUMB_29__14_) );
  FA_X1 u5_mult_82_S2_29_13 ( .A(u5_mult_82_ab_29__13_), .B(
        u5_mult_82_CARRYB_28__13_), .CI(u5_mult_82_SUMB_28__14_), .CO(
        u5_mult_82_CARRYB_29__13_), .S(u5_mult_82_SUMB_29__13_) );
  FA_X1 u5_mult_82_S2_29_12 ( .A(u5_mult_82_ab_29__12_), .B(
        u5_mult_82_CARRYB_28__12_), .CI(u5_mult_82_SUMB_28__13_), .CO(
        u5_mult_82_CARRYB_29__12_), .S(u5_mult_82_SUMB_29__12_) );
  FA_X1 u5_mult_82_S2_29_11 ( .A(u5_mult_82_ab_29__11_), .B(
        u5_mult_82_CARRYB_28__11_), .CI(u5_mult_82_SUMB_28__12_), .CO(
        u5_mult_82_CARRYB_29__11_), .S(u5_mult_82_SUMB_29__11_) );
  FA_X1 u5_mult_82_S2_29_10 ( .A(u5_mult_82_ab_29__10_), .B(
        u5_mult_82_CARRYB_28__10_), .CI(u5_mult_82_SUMB_28__11_), .CO(
        u5_mult_82_CARRYB_29__10_), .S(u5_mult_82_SUMB_29__10_) );
  FA_X1 u5_mult_82_S2_29_9 ( .A(u5_mult_82_ab_29__9_), .B(
        u5_mult_82_CARRYB_28__9_), .CI(u5_mult_82_SUMB_28__10_), .CO(
        u5_mult_82_CARRYB_29__9_), .S(u5_mult_82_SUMB_29__9_) );
  FA_X1 u5_mult_82_S2_29_8 ( .A(u5_mult_82_ab_29__8_), .B(
        u5_mult_82_CARRYB_28__8_), .CI(u5_mult_82_SUMB_28__9_), .CO(
        u5_mult_82_CARRYB_29__8_), .S(u5_mult_82_SUMB_29__8_) );
  FA_X1 u5_mult_82_S2_29_7 ( .A(u5_mult_82_ab_29__7_), .B(
        u5_mult_82_CARRYB_28__7_), .CI(u5_mult_82_SUMB_28__8_), .CO(
        u5_mult_82_CARRYB_29__7_), .S(u5_mult_82_SUMB_29__7_) );
  FA_X1 u5_mult_82_S2_29_6 ( .A(u5_mult_82_ab_29__6_), .B(
        u5_mult_82_CARRYB_28__6_), .CI(u5_mult_82_SUMB_28__7_), .CO(
        u5_mult_82_CARRYB_29__6_), .S(u5_mult_82_SUMB_29__6_) );
  FA_X1 u5_mult_82_S2_29_5 ( .A(u5_mult_82_ab_29__5_), .B(
        u5_mult_82_CARRYB_28__5_), .CI(u5_mult_82_SUMB_28__6_), .CO(
        u5_mult_82_CARRYB_29__5_), .S(u5_mult_82_SUMB_29__5_) );
  FA_X1 u5_mult_82_S2_29_4 ( .A(u5_mult_82_ab_29__4_), .B(
        u5_mult_82_CARRYB_28__4_), .CI(u5_mult_82_SUMB_28__5_), .CO(
        u5_mult_82_CARRYB_29__4_), .S(u5_mult_82_SUMB_29__4_) );
  FA_X1 u5_mult_82_S2_29_3 ( .A(u5_mult_82_ab_29__3_), .B(
        u5_mult_82_CARRYB_28__3_), .CI(u5_mult_82_SUMB_28__4_), .CO(
        u5_mult_82_CARRYB_29__3_), .S(u5_mult_82_SUMB_29__3_) );
  FA_X1 u5_mult_82_S2_29_2 ( .A(u5_mult_82_ab_29__2_), .B(
        u5_mult_82_CARRYB_28__2_), .CI(u5_mult_82_SUMB_28__3_), .CO(
        u5_mult_82_CARRYB_29__2_), .S(u5_mult_82_SUMB_29__2_) );
  FA_X1 u5_mult_82_S2_29_1 ( .A(u5_mult_82_ab_29__1_), .B(
        u5_mult_82_CARRYB_28__1_), .CI(u5_mult_82_SUMB_28__2_), .CO(
        u5_mult_82_CARRYB_29__1_), .S(u5_mult_82_SUMB_29__1_) );
  FA_X1 u5_mult_82_S1_29_0 ( .A(u5_mult_82_ab_29__0_), .B(
        u5_mult_82_CARRYB_28__0_), .CI(u5_mult_82_SUMB_28__1_), .CO(
        u5_mult_82_CARRYB_29__0_), .S(u5_N29) );
  FA_X1 u5_mult_82_S3_30_51 ( .A(u5_mult_82_ab_30__51_), .B(
        u5_mult_82_CARRYB_29__51_), .CI(u5_mult_82_ab_29__52_), .CO(
        u5_mult_82_CARRYB_30__51_), .S(u5_mult_82_SUMB_30__51_) );
  FA_X1 u5_mult_82_S2_30_50 ( .A(u5_mult_82_ab_30__50_), .B(
        u5_mult_82_CARRYB_29__50_), .CI(u5_mult_82_SUMB_29__51_), .CO(
        u5_mult_82_CARRYB_30__50_), .S(u5_mult_82_SUMB_30__50_) );
  FA_X1 u5_mult_82_S2_30_49 ( .A(u5_mult_82_ab_30__49_), .B(
        u5_mult_82_CARRYB_29__49_), .CI(u5_mult_82_SUMB_29__50_), .CO(
        u5_mult_82_CARRYB_30__49_), .S(u5_mult_82_SUMB_30__49_) );
  FA_X1 u5_mult_82_S2_30_48 ( .A(u5_mult_82_ab_30__48_), .B(
        u5_mult_82_CARRYB_29__48_), .CI(u5_mult_82_SUMB_29__49_), .CO(
        u5_mult_82_CARRYB_30__48_), .S(u5_mult_82_SUMB_30__48_) );
  FA_X1 u5_mult_82_S2_30_47 ( .A(u5_mult_82_ab_30__47_), .B(
        u5_mult_82_CARRYB_29__47_), .CI(u5_mult_82_SUMB_29__48_), .CO(
        u5_mult_82_CARRYB_30__47_), .S(u5_mult_82_SUMB_30__47_) );
  FA_X1 u5_mult_82_S2_30_46 ( .A(u5_mult_82_ab_30__46_), .B(
        u5_mult_82_CARRYB_29__46_), .CI(u5_mult_82_SUMB_29__47_), .CO(
        u5_mult_82_CARRYB_30__46_), .S(u5_mult_82_SUMB_30__46_) );
  FA_X1 u5_mult_82_S2_30_45 ( .A(u5_mult_82_ab_30__45_), .B(
        u5_mult_82_CARRYB_29__45_), .CI(u5_mult_82_SUMB_29__46_), .CO(
        u5_mult_82_CARRYB_30__45_), .S(u5_mult_82_SUMB_30__45_) );
  FA_X1 u5_mult_82_S2_30_44 ( .A(u5_mult_82_ab_30__44_), .B(
        u5_mult_82_CARRYB_29__44_), .CI(u5_mult_82_SUMB_29__45_), .CO(
        u5_mult_82_CARRYB_30__44_), .S(u5_mult_82_SUMB_30__44_) );
  FA_X1 u5_mult_82_S2_30_43 ( .A(u5_mult_82_ab_30__43_), .B(
        u5_mult_82_CARRYB_29__43_), .CI(u5_mult_82_SUMB_29__44_), .CO(
        u5_mult_82_CARRYB_30__43_), .S(u5_mult_82_SUMB_30__43_) );
  FA_X1 u5_mult_82_S2_30_42 ( .A(u5_mult_82_ab_30__42_), .B(
        u5_mult_82_CARRYB_29__42_), .CI(u5_mult_82_SUMB_29__43_), .CO(
        u5_mult_82_CARRYB_30__42_), .S(u5_mult_82_SUMB_30__42_) );
  FA_X1 u5_mult_82_S2_30_41 ( .A(u5_mult_82_ab_30__41_), .B(
        u5_mult_82_CARRYB_29__41_), .CI(u5_mult_82_SUMB_29__42_), .CO(
        u5_mult_82_CARRYB_30__41_), .S(u5_mult_82_SUMB_30__41_) );
  FA_X1 u5_mult_82_S2_30_40 ( .A(u5_mult_82_ab_30__40_), .B(
        u5_mult_82_CARRYB_29__40_), .CI(u5_mult_82_SUMB_29__41_), .CO(
        u5_mult_82_CARRYB_30__40_), .S(u5_mult_82_SUMB_30__40_) );
  FA_X1 u5_mult_82_S2_30_39 ( .A(u5_mult_82_ab_30__39_), .B(
        u5_mult_82_CARRYB_29__39_), .CI(u5_mult_82_SUMB_29__40_), .CO(
        u5_mult_82_CARRYB_30__39_), .S(u5_mult_82_SUMB_30__39_) );
  FA_X1 u5_mult_82_S2_30_38 ( .A(u5_mult_82_ab_30__38_), .B(
        u5_mult_82_CARRYB_29__38_), .CI(u5_mult_82_SUMB_29__39_), .CO(
        u5_mult_82_CARRYB_30__38_), .S(u5_mult_82_SUMB_30__38_) );
  FA_X1 u5_mult_82_S2_30_37 ( .A(u5_mult_82_ab_30__37_), .B(
        u5_mult_82_CARRYB_29__37_), .CI(u5_mult_82_SUMB_29__38_), .CO(
        u5_mult_82_CARRYB_30__37_), .S(u5_mult_82_SUMB_30__37_) );
  FA_X1 u5_mult_82_S2_30_36 ( .A(u5_mult_82_ab_30__36_), .B(
        u5_mult_82_CARRYB_29__36_), .CI(u5_mult_82_SUMB_29__37_), .CO(
        u5_mult_82_CARRYB_30__36_), .S(u5_mult_82_SUMB_30__36_) );
  FA_X1 u5_mult_82_S2_30_35 ( .A(u5_mult_82_ab_30__35_), .B(
        u5_mult_82_CARRYB_29__35_), .CI(u5_mult_82_SUMB_29__36_), .CO(
        u5_mult_82_CARRYB_30__35_), .S(u5_mult_82_SUMB_30__35_) );
  FA_X1 u5_mult_82_S2_30_34 ( .A(u5_mult_82_ab_30__34_), .B(
        u5_mult_82_CARRYB_29__34_), .CI(u5_mult_82_SUMB_29__35_), .CO(
        u5_mult_82_CARRYB_30__34_), .S(u5_mult_82_SUMB_30__34_) );
  FA_X1 u5_mult_82_S2_30_33 ( .A(u5_mult_82_ab_30__33_), .B(
        u5_mult_82_CARRYB_29__33_), .CI(u5_mult_82_SUMB_29__34_), .CO(
        u5_mult_82_CARRYB_30__33_), .S(u5_mult_82_SUMB_30__33_) );
  FA_X1 u5_mult_82_S2_30_32 ( .A(u5_mult_82_ab_30__32_), .B(
        u5_mult_82_CARRYB_29__32_), .CI(u5_mult_82_SUMB_29__33_), .CO(
        u5_mult_82_CARRYB_30__32_), .S(u5_mult_82_SUMB_30__32_) );
  FA_X1 u5_mult_82_S2_30_31 ( .A(u5_mult_82_ab_30__31_), .B(
        u5_mult_82_CARRYB_29__31_), .CI(u5_mult_82_SUMB_29__32_), .CO(
        u5_mult_82_CARRYB_30__31_), .S(u5_mult_82_SUMB_30__31_) );
  FA_X1 u5_mult_82_S2_30_30 ( .A(u5_mult_82_ab_30__30_), .B(
        u5_mult_82_CARRYB_29__30_), .CI(u5_mult_82_SUMB_29__31_), .CO(
        u5_mult_82_CARRYB_30__30_), .S(u5_mult_82_SUMB_30__30_) );
  FA_X1 u5_mult_82_S2_30_29 ( .A(u5_mult_82_ab_30__29_), .B(
        u5_mult_82_CARRYB_29__29_), .CI(u5_mult_82_SUMB_29__30_), .CO(
        u5_mult_82_CARRYB_30__29_), .S(u5_mult_82_SUMB_30__29_) );
  FA_X1 u5_mult_82_S2_30_28 ( .A(u5_mult_82_ab_30__28_), .B(
        u5_mult_82_CARRYB_29__28_), .CI(u5_mult_82_SUMB_29__29_), .CO(
        u5_mult_82_CARRYB_30__28_), .S(u5_mult_82_SUMB_30__28_) );
  FA_X1 u5_mult_82_S2_30_27 ( .A(u5_mult_82_ab_30__27_), .B(
        u5_mult_82_CARRYB_29__27_), .CI(u5_mult_82_SUMB_29__28_), .CO(
        u5_mult_82_CARRYB_30__27_), .S(u5_mult_82_SUMB_30__27_) );
  FA_X1 u5_mult_82_S2_30_26 ( .A(u5_mult_82_ab_30__26_), .B(
        u5_mult_82_CARRYB_29__26_), .CI(u5_mult_82_SUMB_29__27_), .CO(
        u5_mult_82_CARRYB_30__26_), .S(u5_mult_82_SUMB_30__26_) );
  FA_X1 u5_mult_82_S2_30_25 ( .A(u5_mult_82_ab_30__25_), .B(
        u5_mult_82_CARRYB_29__25_), .CI(u5_mult_82_SUMB_29__26_), .CO(
        u5_mult_82_CARRYB_30__25_), .S(u5_mult_82_SUMB_30__25_) );
  FA_X1 u5_mult_82_S2_30_24 ( .A(u5_mult_82_ab_30__24_), .B(
        u5_mult_82_CARRYB_29__24_), .CI(u5_mult_82_SUMB_29__25_), .CO(
        u5_mult_82_CARRYB_30__24_), .S(u5_mult_82_SUMB_30__24_) );
  FA_X1 u5_mult_82_S2_30_23 ( .A(u5_mult_82_ab_30__23_), .B(
        u5_mult_82_CARRYB_29__23_), .CI(u5_mult_82_SUMB_29__24_), .CO(
        u5_mult_82_CARRYB_30__23_), .S(u5_mult_82_SUMB_30__23_) );
  FA_X1 u5_mult_82_S2_30_22 ( .A(u5_mult_82_ab_30__22_), .B(
        u5_mult_82_CARRYB_29__22_), .CI(u5_mult_82_SUMB_29__23_), .CO(
        u5_mult_82_CARRYB_30__22_), .S(u5_mult_82_SUMB_30__22_) );
  FA_X1 u5_mult_82_S2_30_21 ( .A(u5_mult_82_ab_30__21_), .B(
        u5_mult_82_CARRYB_29__21_), .CI(u5_mult_82_SUMB_29__22_), .CO(
        u5_mult_82_CARRYB_30__21_), .S(u5_mult_82_SUMB_30__21_) );
  FA_X1 u5_mult_82_S2_30_20 ( .A(u5_mult_82_ab_30__20_), .B(
        u5_mult_82_CARRYB_29__20_), .CI(u5_mult_82_SUMB_29__21_), .CO(
        u5_mult_82_CARRYB_30__20_), .S(u5_mult_82_SUMB_30__20_) );
  FA_X1 u5_mult_82_S2_30_19 ( .A(u5_mult_82_ab_30__19_), .B(
        u5_mult_82_CARRYB_29__19_), .CI(u5_mult_82_SUMB_29__20_), .CO(
        u5_mult_82_CARRYB_30__19_), .S(u5_mult_82_SUMB_30__19_) );
  FA_X1 u5_mult_82_S2_30_18 ( .A(u5_mult_82_ab_30__18_), .B(
        u5_mult_82_CARRYB_29__18_), .CI(u5_mult_82_SUMB_29__19_), .CO(
        u5_mult_82_CARRYB_30__18_), .S(u5_mult_82_SUMB_30__18_) );
  FA_X1 u5_mult_82_S2_30_17 ( .A(u5_mult_82_ab_30__17_), .B(
        u5_mult_82_CARRYB_29__17_), .CI(u5_mult_82_SUMB_29__18_), .CO(
        u5_mult_82_CARRYB_30__17_), .S(u5_mult_82_SUMB_30__17_) );
  FA_X1 u5_mult_82_S2_30_16 ( .A(u5_mult_82_ab_30__16_), .B(
        u5_mult_82_CARRYB_29__16_), .CI(u5_mult_82_SUMB_29__17_), .CO(
        u5_mult_82_CARRYB_30__16_), .S(u5_mult_82_SUMB_30__16_) );
  FA_X1 u5_mult_82_S2_30_15 ( .A(u5_mult_82_ab_30__15_), .B(
        u5_mult_82_CARRYB_29__15_), .CI(u5_mult_82_SUMB_29__16_), .CO(
        u5_mult_82_CARRYB_30__15_), .S(u5_mult_82_SUMB_30__15_) );
  FA_X1 u5_mult_82_S2_30_14 ( .A(u5_mult_82_ab_30__14_), .B(
        u5_mult_82_CARRYB_29__14_), .CI(u5_mult_82_SUMB_29__15_), .CO(
        u5_mult_82_CARRYB_30__14_), .S(u5_mult_82_SUMB_30__14_) );
  FA_X1 u5_mult_82_S2_30_13 ( .A(u5_mult_82_ab_30__13_), .B(
        u5_mult_82_CARRYB_29__13_), .CI(u5_mult_82_SUMB_29__14_), .CO(
        u5_mult_82_CARRYB_30__13_), .S(u5_mult_82_SUMB_30__13_) );
  FA_X1 u5_mult_82_S2_30_12 ( .A(u5_mult_82_ab_30__12_), .B(
        u5_mult_82_CARRYB_29__12_), .CI(u5_mult_82_SUMB_29__13_), .CO(
        u5_mult_82_CARRYB_30__12_), .S(u5_mult_82_SUMB_30__12_) );
  FA_X1 u5_mult_82_S2_30_11 ( .A(u5_mult_82_ab_30__11_), .B(
        u5_mult_82_CARRYB_29__11_), .CI(u5_mult_82_SUMB_29__12_), .CO(
        u5_mult_82_CARRYB_30__11_), .S(u5_mult_82_SUMB_30__11_) );
  FA_X1 u5_mult_82_S2_30_10 ( .A(u5_mult_82_ab_30__10_), .B(
        u5_mult_82_CARRYB_29__10_), .CI(u5_mult_82_SUMB_29__11_), .CO(
        u5_mult_82_CARRYB_30__10_), .S(u5_mult_82_SUMB_30__10_) );
  FA_X1 u5_mult_82_S2_30_9 ( .A(u5_mult_82_ab_30__9_), .B(
        u5_mult_82_CARRYB_29__9_), .CI(u5_mult_82_SUMB_29__10_), .CO(
        u5_mult_82_CARRYB_30__9_), .S(u5_mult_82_SUMB_30__9_) );
  FA_X1 u5_mult_82_S2_30_8 ( .A(u5_mult_82_ab_30__8_), .B(
        u5_mult_82_CARRYB_29__8_), .CI(u5_mult_82_SUMB_29__9_), .CO(
        u5_mult_82_CARRYB_30__8_), .S(u5_mult_82_SUMB_30__8_) );
  FA_X1 u5_mult_82_S2_30_7 ( .A(u5_mult_82_ab_30__7_), .B(
        u5_mult_82_CARRYB_29__7_), .CI(u5_mult_82_SUMB_29__8_), .CO(
        u5_mult_82_CARRYB_30__7_), .S(u5_mult_82_SUMB_30__7_) );
  FA_X1 u5_mult_82_S2_30_6 ( .A(u5_mult_82_ab_30__6_), .B(
        u5_mult_82_CARRYB_29__6_), .CI(u5_mult_82_SUMB_29__7_), .CO(
        u5_mult_82_CARRYB_30__6_), .S(u5_mult_82_SUMB_30__6_) );
  FA_X1 u5_mult_82_S2_30_5 ( .A(u5_mult_82_ab_30__5_), .B(
        u5_mult_82_CARRYB_29__5_), .CI(u5_mult_82_SUMB_29__6_), .CO(
        u5_mult_82_CARRYB_30__5_), .S(u5_mult_82_SUMB_30__5_) );
  FA_X1 u5_mult_82_S2_30_4 ( .A(u5_mult_82_ab_30__4_), .B(
        u5_mult_82_CARRYB_29__4_), .CI(u5_mult_82_SUMB_29__5_), .CO(
        u5_mult_82_CARRYB_30__4_), .S(u5_mult_82_SUMB_30__4_) );
  FA_X1 u5_mult_82_S2_30_3 ( .A(u5_mult_82_ab_30__3_), .B(
        u5_mult_82_CARRYB_29__3_), .CI(u5_mult_82_SUMB_29__4_), .CO(
        u5_mult_82_CARRYB_30__3_), .S(u5_mult_82_SUMB_30__3_) );
  FA_X1 u5_mult_82_S2_30_2 ( .A(u5_mult_82_ab_30__2_), .B(
        u5_mult_82_CARRYB_29__2_), .CI(u5_mult_82_SUMB_29__3_), .CO(
        u5_mult_82_CARRYB_30__2_), .S(u5_mult_82_SUMB_30__2_) );
  FA_X1 u5_mult_82_S2_30_1 ( .A(u5_mult_82_ab_30__1_), .B(
        u5_mult_82_CARRYB_29__1_), .CI(u5_mult_82_SUMB_29__2_), .CO(
        u5_mult_82_CARRYB_30__1_), .S(u5_mult_82_SUMB_30__1_) );
  FA_X1 u5_mult_82_S1_30_0 ( .A(u5_mult_82_ab_30__0_), .B(
        u5_mult_82_CARRYB_29__0_), .CI(u5_mult_82_SUMB_29__1_), .CO(
        u5_mult_82_CARRYB_30__0_), .S(u5_N30) );
  FA_X1 u5_mult_82_S3_31_51 ( .A(u5_mult_82_ab_31__51_), .B(
        u5_mult_82_CARRYB_30__51_), .CI(u5_mult_82_ab_30__52_), .CO(
        u5_mult_82_CARRYB_31__51_), .S(u5_mult_82_SUMB_31__51_) );
  FA_X1 u5_mult_82_S2_31_50 ( .A(u5_mult_82_ab_31__50_), .B(
        u5_mult_82_CARRYB_30__50_), .CI(u5_mult_82_SUMB_30__51_), .CO(
        u5_mult_82_CARRYB_31__50_), .S(u5_mult_82_SUMB_31__50_) );
  FA_X1 u5_mult_82_S2_31_49 ( .A(u5_mult_82_ab_31__49_), .B(
        u5_mult_82_CARRYB_30__49_), .CI(u5_mult_82_SUMB_30__50_), .CO(
        u5_mult_82_CARRYB_31__49_), .S(u5_mult_82_SUMB_31__49_) );
  FA_X1 u5_mult_82_S2_31_48 ( .A(u5_mult_82_ab_31__48_), .B(
        u5_mult_82_CARRYB_30__48_), .CI(u5_mult_82_SUMB_30__49_), .CO(
        u5_mult_82_CARRYB_31__48_), .S(u5_mult_82_SUMB_31__48_) );
  FA_X1 u5_mult_82_S2_31_47 ( .A(u5_mult_82_ab_31__47_), .B(
        u5_mult_82_CARRYB_30__47_), .CI(u5_mult_82_SUMB_30__48_), .CO(
        u5_mult_82_CARRYB_31__47_), .S(u5_mult_82_SUMB_31__47_) );
  FA_X1 u5_mult_82_S2_31_46 ( .A(u5_mult_82_ab_31__46_), .B(
        u5_mult_82_CARRYB_30__46_), .CI(u5_mult_82_SUMB_30__47_), .CO(
        u5_mult_82_CARRYB_31__46_), .S(u5_mult_82_SUMB_31__46_) );
  FA_X1 u5_mult_82_S2_31_45 ( .A(u5_mult_82_ab_31__45_), .B(
        u5_mult_82_CARRYB_30__45_), .CI(u5_mult_82_SUMB_30__46_), .CO(
        u5_mult_82_CARRYB_31__45_), .S(u5_mult_82_SUMB_31__45_) );
  FA_X1 u5_mult_82_S2_31_44 ( .A(u5_mult_82_ab_31__44_), .B(
        u5_mult_82_CARRYB_30__44_), .CI(u5_mult_82_SUMB_30__45_), .CO(
        u5_mult_82_CARRYB_31__44_), .S(u5_mult_82_SUMB_31__44_) );
  FA_X1 u5_mult_82_S2_31_43 ( .A(u5_mult_82_ab_31__43_), .B(
        u5_mult_82_CARRYB_30__43_), .CI(u5_mult_82_SUMB_30__44_), .CO(
        u5_mult_82_CARRYB_31__43_), .S(u5_mult_82_SUMB_31__43_) );
  FA_X1 u5_mult_82_S2_31_42 ( .A(u5_mult_82_ab_31__42_), .B(
        u5_mult_82_CARRYB_30__42_), .CI(u5_mult_82_SUMB_30__43_), .CO(
        u5_mult_82_CARRYB_31__42_), .S(u5_mult_82_SUMB_31__42_) );
  FA_X1 u5_mult_82_S2_31_41 ( .A(u5_mult_82_ab_31__41_), .B(
        u5_mult_82_CARRYB_30__41_), .CI(u5_mult_82_SUMB_30__42_), .CO(
        u5_mult_82_CARRYB_31__41_), .S(u5_mult_82_SUMB_31__41_) );
  FA_X1 u5_mult_82_S2_31_40 ( .A(u5_mult_82_ab_31__40_), .B(
        u5_mult_82_CARRYB_30__40_), .CI(u5_mult_82_SUMB_30__41_), .CO(
        u5_mult_82_CARRYB_31__40_), .S(u5_mult_82_SUMB_31__40_) );
  FA_X1 u5_mult_82_S2_31_39 ( .A(u5_mult_82_ab_31__39_), .B(
        u5_mult_82_CARRYB_30__39_), .CI(u5_mult_82_SUMB_30__40_), .CO(
        u5_mult_82_CARRYB_31__39_), .S(u5_mult_82_SUMB_31__39_) );
  FA_X1 u5_mult_82_S2_31_38 ( .A(u5_mult_82_ab_31__38_), .B(
        u5_mult_82_CARRYB_30__38_), .CI(u5_mult_82_SUMB_30__39_), .CO(
        u5_mult_82_CARRYB_31__38_), .S(u5_mult_82_SUMB_31__38_) );
  FA_X1 u5_mult_82_S2_31_37 ( .A(u5_mult_82_ab_31__37_), .B(
        u5_mult_82_CARRYB_30__37_), .CI(u5_mult_82_SUMB_30__38_), .CO(
        u5_mult_82_CARRYB_31__37_), .S(u5_mult_82_SUMB_31__37_) );
  FA_X1 u5_mult_82_S2_31_36 ( .A(u5_mult_82_ab_31__36_), .B(
        u5_mult_82_CARRYB_30__36_), .CI(u5_mult_82_SUMB_30__37_), .CO(
        u5_mult_82_CARRYB_31__36_), .S(u5_mult_82_SUMB_31__36_) );
  FA_X1 u5_mult_82_S2_31_35 ( .A(u5_mult_82_ab_31__35_), .B(
        u5_mult_82_CARRYB_30__35_), .CI(u5_mult_82_SUMB_30__36_), .CO(
        u5_mult_82_CARRYB_31__35_), .S(u5_mult_82_SUMB_31__35_) );
  FA_X1 u5_mult_82_S2_31_34 ( .A(u5_mult_82_ab_31__34_), .B(
        u5_mult_82_CARRYB_30__34_), .CI(u5_mult_82_SUMB_30__35_), .CO(
        u5_mult_82_CARRYB_31__34_), .S(u5_mult_82_SUMB_31__34_) );
  FA_X1 u5_mult_82_S2_31_33 ( .A(u5_mult_82_ab_31__33_), .B(
        u5_mult_82_CARRYB_30__33_), .CI(u5_mult_82_SUMB_30__34_), .CO(
        u5_mult_82_CARRYB_31__33_), .S(u5_mult_82_SUMB_31__33_) );
  FA_X1 u5_mult_82_S2_31_32 ( .A(u5_mult_82_ab_31__32_), .B(
        u5_mult_82_CARRYB_30__32_), .CI(u5_mult_82_SUMB_30__33_), .CO(
        u5_mult_82_CARRYB_31__32_), .S(u5_mult_82_SUMB_31__32_) );
  FA_X1 u5_mult_82_S2_31_31 ( .A(u5_mult_82_ab_31__31_), .B(
        u5_mult_82_CARRYB_30__31_), .CI(u5_mult_82_SUMB_30__32_), .CO(
        u5_mult_82_CARRYB_31__31_), .S(u5_mult_82_SUMB_31__31_) );
  FA_X1 u5_mult_82_S2_31_30 ( .A(u5_mult_82_ab_31__30_), .B(
        u5_mult_82_CARRYB_30__30_), .CI(u5_mult_82_SUMB_30__31_), .CO(
        u5_mult_82_CARRYB_31__30_), .S(u5_mult_82_SUMB_31__30_) );
  FA_X1 u5_mult_82_S2_31_29 ( .A(u5_mult_82_ab_31__29_), .B(
        u5_mult_82_CARRYB_30__29_), .CI(u5_mult_82_SUMB_30__30_), .CO(
        u5_mult_82_CARRYB_31__29_), .S(u5_mult_82_SUMB_31__29_) );
  FA_X1 u5_mult_82_S2_31_28 ( .A(u5_mult_82_ab_31__28_), .B(
        u5_mult_82_CARRYB_30__28_), .CI(u5_mult_82_SUMB_30__29_), .CO(
        u5_mult_82_CARRYB_31__28_), .S(u5_mult_82_SUMB_31__28_) );
  FA_X1 u5_mult_82_S2_31_27 ( .A(u5_mult_82_ab_31__27_), .B(
        u5_mult_82_CARRYB_30__27_), .CI(u5_mult_82_SUMB_30__28_), .CO(
        u5_mult_82_CARRYB_31__27_), .S(u5_mult_82_SUMB_31__27_) );
  FA_X1 u5_mult_82_S2_31_26 ( .A(u5_mult_82_ab_31__26_), .B(
        u5_mult_82_CARRYB_30__26_), .CI(u5_mult_82_SUMB_30__27_), .CO(
        u5_mult_82_CARRYB_31__26_), .S(u5_mult_82_SUMB_31__26_) );
  FA_X1 u5_mult_82_S2_31_25 ( .A(u5_mult_82_ab_31__25_), .B(
        u5_mult_82_CARRYB_30__25_), .CI(u5_mult_82_SUMB_30__26_), .CO(
        u5_mult_82_CARRYB_31__25_), .S(u5_mult_82_SUMB_31__25_) );
  FA_X1 u5_mult_82_S2_31_24 ( .A(u5_mult_82_ab_31__24_), .B(
        u5_mult_82_CARRYB_30__24_), .CI(u5_mult_82_SUMB_30__25_), .CO(
        u5_mult_82_CARRYB_31__24_), .S(u5_mult_82_SUMB_31__24_) );
  FA_X1 u5_mult_82_S2_31_23 ( .A(u5_mult_82_ab_31__23_), .B(
        u5_mult_82_CARRYB_30__23_), .CI(u5_mult_82_SUMB_30__24_), .CO(
        u5_mult_82_CARRYB_31__23_), .S(u5_mult_82_SUMB_31__23_) );
  FA_X1 u5_mult_82_S2_31_22 ( .A(u5_mult_82_ab_31__22_), .B(
        u5_mult_82_CARRYB_30__22_), .CI(u5_mult_82_SUMB_30__23_), .CO(
        u5_mult_82_CARRYB_31__22_), .S(u5_mult_82_SUMB_31__22_) );
  FA_X1 u5_mult_82_S2_31_21 ( .A(u5_mult_82_ab_31__21_), .B(
        u5_mult_82_CARRYB_30__21_), .CI(u5_mult_82_SUMB_30__22_), .CO(
        u5_mult_82_CARRYB_31__21_), .S(u5_mult_82_SUMB_31__21_) );
  FA_X1 u5_mult_82_S2_31_20 ( .A(u5_mult_82_ab_31__20_), .B(
        u5_mult_82_CARRYB_30__20_), .CI(u5_mult_82_SUMB_30__21_), .CO(
        u5_mult_82_CARRYB_31__20_), .S(u5_mult_82_SUMB_31__20_) );
  FA_X1 u5_mult_82_S2_31_19 ( .A(u5_mult_82_ab_31__19_), .B(
        u5_mult_82_CARRYB_30__19_), .CI(u5_mult_82_SUMB_30__20_), .CO(
        u5_mult_82_CARRYB_31__19_), .S(u5_mult_82_SUMB_31__19_) );
  FA_X1 u5_mult_82_S2_31_18 ( .A(u5_mult_82_ab_31__18_), .B(
        u5_mult_82_CARRYB_30__18_), .CI(u5_mult_82_SUMB_30__19_), .CO(
        u5_mult_82_CARRYB_31__18_), .S(u5_mult_82_SUMB_31__18_) );
  FA_X1 u5_mult_82_S2_31_17 ( .A(u5_mult_82_ab_31__17_), .B(
        u5_mult_82_CARRYB_30__17_), .CI(u5_mult_82_SUMB_30__18_), .CO(
        u5_mult_82_CARRYB_31__17_), .S(u5_mult_82_SUMB_31__17_) );
  FA_X1 u5_mult_82_S2_31_16 ( .A(u5_mult_82_ab_31__16_), .B(
        u5_mult_82_CARRYB_30__16_), .CI(u5_mult_82_SUMB_30__17_), .CO(
        u5_mult_82_CARRYB_31__16_), .S(u5_mult_82_SUMB_31__16_) );
  FA_X1 u5_mult_82_S2_31_15 ( .A(u5_mult_82_ab_31__15_), .B(
        u5_mult_82_CARRYB_30__15_), .CI(u5_mult_82_SUMB_30__16_), .CO(
        u5_mult_82_CARRYB_31__15_), .S(u5_mult_82_SUMB_31__15_) );
  FA_X1 u5_mult_82_S2_31_14 ( .A(u5_mult_82_ab_31__14_), .B(
        u5_mult_82_CARRYB_30__14_), .CI(u5_mult_82_SUMB_30__15_), .CO(
        u5_mult_82_CARRYB_31__14_), .S(u5_mult_82_SUMB_31__14_) );
  FA_X1 u5_mult_82_S2_31_13 ( .A(u5_mult_82_ab_31__13_), .B(
        u5_mult_82_CARRYB_30__13_), .CI(u5_mult_82_SUMB_30__14_), .CO(
        u5_mult_82_CARRYB_31__13_), .S(u5_mult_82_SUMB_31__13_) );
  FA_X1 u5_mult_82_S2_31_12 ( .A(u5_mult_82_ab_31__12_), .B(
        u5_mult_82_CARRYB_30__12_), .CI(u5_mult_82_SUMB_30__13_), .CO(
        u5_mult_82_CARRYB_31__12_), .S(u5_mult_82_SUMB_31__12_) );
  FA_X1 u5_mult_82_S2_31_11 ( .A(u5_mult_82_ab_31__11_), .B(
        u5_mult_82_CARRYB_30__11_), .CI(u5_mult_82_SUMB_30__12_), .CO(
        u5_mult_82_CARRYB_31__11_), .S(u5_mult_82_SUMB_31__11_) );
  FA_X1 u5_mult_82_S2_31_10 ( .A(u5_mult_82_ab_31__10_), .B(
        u5_mult_82_CARRYB_30__10_), .CI(u5_mult_82_SUMB_30__11_), .CO(
        u5_mult_82_CARRYB_31__10_), .S(u5_mult_82_SUMB_31__10_) );
  FA_X1 u5_mult_82_S2_31_9 ( .A(u5_mult_82_ab_31__9_), .B(
        u5_mult_82_CARRYB_30__9_), .CI(u5_mult_82_SUMB_30__10_), .CO(
        u5_mult_82_CARRYB_31__9_), .S(u5_mult_82_SUMB_31__9_) );
  FA_X1 u5_mult_82_S2_31_8 ( .A(u5_mult_82_ab_31__8_), .B(
        u5_mult_82_CARRYB_30__8_), .CI(u5_mult_82_SUMB_30__9_), .CO(
        u5_mult_82_CARRYB_31__8_), .S(u5_mult_82_SUMB_31__8_) );
  FA_X1 u5_mult_82_S2_31_7 ( .A(u5_mult_82_ab_31__7_), .B(
        u5_mult_82_CARRYB_30__7_), .CI(u5_mult_82_SUMB_30__8_), .CO(
        u5_mult_82_CARRYB_31__7_), .S(u5_mult_82_SUMB_31__7_) );
  FA_X1 u5_mult_82_S2_31_6 ( .A(u5_mult_82_ab_31__6_), .B(
        u5_mult_82_CARRYB_30__6_), .CI(u5_mult_82_SUMB_30__7_), .CO(
        u5_mult_82_CARRYB_31__6_), .S(u5_mult_82_SUMB_31__6_) );
  FA_X1 u5_mult_82_S2_31_5 ( .A(u5_mult_82_ab_31__5_), .B(
        u5_mult_82_CARRYB_30__5_), .CI(u5_mult_82_SUMB_30__6_), .CO(
        u5_mult_82_CARRYB_31__5_), .S(u5_mult_82_SUMB_31__5_) );
  FA_X1 u5_mult_82_S2_31_4 ( .A(u5_mult_82_ab_31__4_), .B(
        u5_mult_82_CARRYB_30__4_), .CI(u5_mult_82_SUMB_30__5_), .CO(
        u5_mult_82_CARRYB_31__4_), .S(u5_mult_82_SUMB_31__4_) );
  FA_X1 u5_mult_82_S2_31_3 ( .A(u5_mult_82_ab_31__3_), .B(
        u5_mult_82_CARRYB_30__3_), .CI(u5_mult_82_SUMB_30__4_), .CO(
        u5_mult_82_CARRYB_31__3_), .S(u5_mult_82_SUMB_31__3_) );
  FA_X1 u5_mult_82_S2_31_2 ( .A(u5_mult_82_ab_31__2_), .B(
        u5_mult_82_CARRYB_30__2_), .CI(u5_mult_82_SUMB_30__3_), .CO(
        u5_mult_82_CARRYB_31__2_), .S(u5_mult_82_SUMB_31__2_) );
  FA_X1 u5_mult_82_S2_31_1 ( .A(u5_mult_82_ab_31__1_), .B(
        u5_mult_82_CARRYB_30__1_), .CI(u5_mult_82_SUMB_30__2_), .CO(
        u5_mult_82_CARRYB_31__1_), .S(u5_mult_82_SUMB_31__1_) );
  FA_X1 u5_mult_82_S1_31_0 ( .A(u5_mult_82_ab_31__0_), .B(
        u5_mult_82_CARRYB_30__0_), .CI(u5_mult_82_SUMB_30__1_), .CO(
        u5_mult_82_CARRYB_31__0_), .S(u5_N31) );
  FA_X1 u5_mult_82_S3_32_51 ( .A(u5_mult_82_ab_32__51_), .B(
        u5_mult_82_CARRYB_31__51_), .CI(u5_mult_82_ab_31__52_), .CO(
        u5_mult_82_CARRYB_32__51_), .S(u5_mult_82_SUMB_32__51_) );
  FA_X1 u5_mult_82_S2_32_50 ( .A(u5_mult_82_ab_32__50_), .B(
        u5_mult_82_CARRYB_31__50_), .CI(u5_mult_82_SUMB_31__51_), .CO(
        u5_mult_82_CARRYB_32__50_), .S(u5_mult_82_SUMB_32__50_) );
  FA_X1 u5_mult_82_S2_32_49 ( .A(u5_mult_82_ab_32__49_), .B(
        u5_mult_82_CARRYB_31__49_), .CI(u5_mult_82_SUMB_31__50_), .CO(
        u5_mult_82_CARRYB_32__49_), .S(u5_mult_82_SUMB_32__49_) );
  FA_X1 u5_mult_82_S2_32_48 ( .A(u5_mult_82_ab_32__48_), .B(
        u5_mult_82_CARRYB_31__48_), .CI(u5_mult_82_SUMB_31__49_), .CO(
        u5_mult_82_CARRYB_32__48_), .S(u5_mult_82_SUMB_32__48_) );
  FA_X1 u5_mult_82_S2_32_47 ( .A(u5_mult_82_ab_32__47_), .B(
        u5_mult_82_CARRYB_31__47_), .CI(u5_mult_82_SUMB_31__48_), .CO(
        u5_mult_82_CARRYB_32__47_), .S(u5_mult_82_SUMB_32__47_) );
  FA_X1 u5_mult_82_S2_32_46 ( .A(u5_mult_82_ab_32__46_), .B(
        u5_mult_82_CARRYB_31__46_), .CI(u5_mult_82_SUMB_31__47_), .CO(
        u5_mult_82_CARRYB_32__46_), .S(u5_mult_82_SUMB_32__46_) );
  FA_X1 u5_mult_82_S2_32_45 ( .A(u5_mult_82_ab_32__45_), .B(
        u5_mult_82_CARRYB_31__45_), .CI(u5_mult_82_SUMB_31__46_), .CO(
        u5_mult_82_CARRYB_32__45_), .S(u5_mult_82_SUMB_32__45_) );
  FA_X1 u5_mult_82_S2_32_44 ( .A(u5_mult_82_ab_32__44_), .B(
        u5_mult_82_CARRYB_31__44_), .CI(u5_mult_82_SUMB_31__45_), .CO(
        u5_mult_82_CARRYB_32__44_), .S(u5_mult_82_SUMB_32__44_) );
  FA_X1 u5_mult_82_S2_32_43 ( .A(u5_mult_82_ab_32__43_), .B(
        u5_mult_82_CARRYB_31__43_), .CI(u5_mult_82_SUMB_31__44_), .CO(
        u5_mult_82_CARRYB_32__43_), .S(u5_mult_82_SUMB_32__43_) );
  FA_X1 u5_mult_82_S2_32_42 ( .A(u5_mult_82_ab_32__42_), .B(
        u5_mult_82_CARRYB_31__42_), .CI(u5_mult_82_SUMB_31__43_), .CO(
        u5_mult_82_CARRYB_32__42_), .S(u5_mult_82_SUMB_32__42_) );
  FA_X1 u5_mult_82_S2_32_41 ( .A(u5_mult_82_ab_32__41_), .B(
        u5_mult_82_CARRYB_31__41_), .CI(u5_mult_82_SUMB_31__42_), .CO(
        u5_mult_82_CARRYB_32__41_), .S(u5_mult_82_SUMB_32__41_) );
  FA_X1 u5_mult_82_S2_32_40 ( .A(u5_mult_82_ab_32__40_), .B(
        u5_mult_82_CARRYB_31__40_), .CI(u5_mult_82_SUMB_31__41_), .CO(
        u5_mult_82_CARRYB_32__40_), .S(u5_mult_82_SUMB_32__40_) );
  FA_X1 u5_mult_82_S2_32_39 ( .A(u5_mult_82_ab_32__39_), .B(
        u5_mult_82_CARRYB_31__39_), .CI(u5_mult_82_SUMB_31__40_), .CO(
        u5_mult_82_CARRYB_32__39_), .S(u5_mult_82_SUMB_32__39_) );
  FA_X1 u5_mult_82_S2_32_38 ( .A(u5_mult_82_ab_32__38_), .B(
        u5_mult_82_CARRYB_31__38_), .CI(u5_mult_82_SUMB_31__39_), .CO(
        u5_mult_82_CARRYB_32__38_), .S(u5_mult_82_SUMB_32__38_) );
  FA_X1 u5_mult_82_S2_32_37 ( .A(u5_mult_82_ab_32__37_), .B(
        u5_mult_82_CARRYB_31__37_), .CI(u5_mult_82_SUMB_31__38_), .CO(
        u5_mult_82_CARRYB_32__37_), .S(u5_mult_82_SUMB_32__37_) );
  FA_X1 u5_mult_82_S2_32_36 ( .A(u5_mult_82_ab_32__36_), .B(
        u5_mult_82_CARRYB_31__36_), .CI(u5_mult_82_SUMB_31__37_), .CO(
        u5_mult_82_CARRYB_32__36_), .S(u5_mult_82_SUMB_32__36_) );
  FA_X1 u5_mult_82_S2_32_35 ( .A(u5_mult_82_ab_32__35_), .B(
        u5_mult_82_CARRYB_31__35_), .CI(u5_mult_82_SUMB_31__36_), .CO(
        u5_mult_82_CARRYB_32__35_), .S(u5_mult_82_SUMB_32__35_) );
  FA_X1 u5_mult_82_S2_32_34 ( .A(u5_mult_82_ab_32__34_), .B(
        u5_mult_82_CARRYB_31__34_), .CI(u5_mult_82_SUMB_31__35_), .CO(
        u5_mult_82_CARRYB_32__34_), .S(u5_mult_82_SUMB_32__34_) );
  FA_X1 u5_mult_82_S2_32_33 ( .A(u5_mult_82_ab_32__33_), .B(
        u5_mult_82_CARRYB_31__33_), .CI(u5_mult_82_SUMB_31__34_), .CO(
        u5_mult_82_CARRYB_32__33_), .S(u5_mult_82_SUMB_32__33_) );
  FA_X1 u5_mult_82_S2_32_32 ( .A(u5_mult_82_ab_32__32_), .B(
        u5_mult_82_CARRYB_31__32_), .CI(u5_mult_82_SUMB_31__33_), .CO(
        u5_mult_82_CARRYB_32__32_), .S(u5_mult_82_SUMB_32__32_) );
  FA_X1 u5_mult_82_S2_32_31 ( .A(u5_mult_82_ab_32__31_), .B(
        u5_mult_82_CARRYB_31__31_), .CI(u5_mult_82_SUMB_31__32_), .CO(
        u5_mult_82_CARRYB_32__31_), .S(u5_mult_82_SUMB_32__31_) );
  FA_X1 u5_mult_82_S2_32_30 ( .A(u5_mult_82_ab_32__30_), .B(
        u5_mult_82_CARRYB_31__30_), .CI(u5_mult_82_SUMB_31__31_), .CO(
        u5_mult_82_CARRYB_32__30_), .S(u5_mult_82_SUMB_32__30_) );
  FA_X1 u5_mult_82_S2_32_29 ( .A(u5_mult_82_ab_32__29_), .B(
        u5_mult_82_CARRYB_31__29_), .CI(u5_mult_82_SUMB_31__30_), .CO(
        u5_mult_82_CARRYB_32__29_), .S(u5_mult_82_SUMB_32__29_) );
  FA_X1 u5_mult_82_S2_32_28 ( .A(u5_mult_82_ab_32__28_), .B(
        u5_mult_82_CARRYB_31__28_), .CI(u5_mult_82_SUMB_31__29_), .CO(
        u5_mult_82_CARRYB_32__28_), .S(u5_mult_82_SUMB_32__28_) );
  FA_X1 u5_mult_82_S2_32_27 ( .A(u5_mult_82_ab_32__27_), .B(
        u5_mult_82_CARRYB_31__27_), .CI(u5_mult_82_SUMB_31__28_), .CO(
        u5_mult_82_CARRYB_32__27_), .S(u5_mult_82_SUMB_32__27_) );
  FA_X1 u5_mult_82_S2_32_26 ( .A(u5_mult_82_ab_32__26_), .B(
        u5_mult_82_CARRYB_31__26_), .CI(u5_mult_82_SUMB_31__27_), .CO(
        u5_mult_82_CARRYB_32__26_), .S(u5_mult_82_SUMB_32__26_) );
  FA_X1 u5_mult_82_S2_32_25 ( .A(u5_mult_82_ab_32__25_), .B(
        u5_mult_82_CARRYB_31__25_), .CI(u5_mult_82_SUMB_31__26_), .CO(
        u5_mult_82_CARRYB_32__25_), .S(u5_mult_82_SUMB_32__25_) );
  FA_X1 u5_mult_82_S2_32_24 ( .A(u5_mult_82_ab_32__24_), .B(
        u5_mult_82_CARRYB_31__24_), .CI(u5_mult_82_SUMB_31__25_), .CO(
        u5_mult_82_CARRYB_32__24_), .S(u5_mult_82_SUMB_32__24_) );
  FA_X1 u5_mult_82_S2_32_23 ( .A(u5_mult_82_ab_32__23_), .B(
        u5_mult_82_CARRYB_31__23_), .CI(u5_mult_82_SUMB_31__24_), .CO(
        u5_mult_82_CARRYB_32__23_), .S(u5_mult_82_SUMB_32__23_) );
  FA_X1 u5_mult_82_S2_32_22 ( .A(u5_mult_82_ab_32__22_), .B(
        u5_mult_82_CARRYB_31__22_), .CI(u5_mult_82_SUMB_31__23_), .CO(
        u5_mult_82_CARRYB_32__22_), .S(u5_mult_82_SUMB_32__22_) );
  FA_X1 u5_mult_82_S2_32_21 ( .A(u5_mult_82_ab_32__21_), .B(
        u5_mult_82_CARRYB_31__21_), .CI(u5_mult_82_SUMB_31__22_), .CO(
        u5_mult_82_CARRYB_32__21_), .S(u5_mult_82_SUMB_32__21_) );
  FA_X1 u5_mult_82_S2_32_20 ( .A(u5_mult_82_ab_32__20_), .B(
        u5_mult_82_CARRYB_31__20_), .CI(u5_mult_82_SUMB_31__21_), .CO(
        u5_mult_82_CARRYB_32__20_), .S(u5_mult_82_SUMB_32__20_) );
  FA_X1 u5_mult_82_S2_32_19 ( .A(u5_mult_82_ab_32__19_), .B(
        u5_mult_82_CARRYB_31__19_), .CI(u5_mult_82_SUMB_31__20_), .CO(
        u5_mult_82_CARRYB_32__19_), .S(u5_mult_82_SUMB_32__19_) );
  FA_X1 u5_mult_82_S2_32_18 ( .A(u5_mult_82_ab_32__18_), .B(
        u5_mult_82_CARRYB_31__18_), .CI(u5_mult_82_SUMB_31__19_), .CO(
        u5_mult_82_CARRYB_32__18_), .S(u5_mult_82_SUMB_32__18_) );
  FA_X1 u5_mult_82_S2_32_17 ( .A(u5_mult_82_ab_32__17_), .B(
        u5_mult_82_CARRYB_31__17_), .CI(u5_mult_82_SUMB_31__18_), .CO(
        u5_mult_82_CARRYB_32__17_), .S(u5_mult_82_SUMB_32__17_) );
  FA_X1 u5_mult_82_S2_32_16 ( .A(u5_mult_82_ab_32__16_), .B(
        u5_mult_82_CARRYB_31__16_), .CI(u5_mult_82_SUMB_31__17_), .CO(
        u5_mult_82_CARRYB_32__16_), .S(u5_mult_82_SUMB_32__16_) );
  FA_X1 u5_mult_82_S2_32_15 ( .A(u5_mult_82_ab_32__15_), .B(
        u5_mult_82_CARRYB_31__15_), .CI(u5_mult_82_SUMB_31__16_), .CO(
        u5_mult_82_CARRYB_32__15_), .S(u5_mult_82_SUMB_32__15_) );
  FA_X1 u5_mult_82_S2_32_14 ( .A(u5_mult_82_ab_32__14_), .B(
        u5_mult_82_CARRYB_31__14_), .CI(u5_mult_82_SUMB_31__15_), .CO(
        u5_mult_82_CARRYB_32__14_), .S(u5_mult_82_SUMB_32__14_) );
  FA_X1 u5_mult_82_S2_32_13 ( .A(u5_mult_82_ab_32__13_), .B(
        u5_mult_82_CARRYB_31__13_), .CI(u5_mult_82_SUMB_31__14_), .CO(
        u5_mult_82_CARRYB_32__13_), .S(u5_mult_82_SUMB_32__13_) );
  FA_X1 u5_mult_82_S2_32_12 ( .A(u5_mult_82_ab_32__12_), .B(
        u5_mult_82_CARRYB_31__12_), .CI(u5_mult_82_SUMB_31__13_), .CO(
        u5_mult_82_CARRYB_32__12_), .S(u5_mult_82_SUMB_32__12_) );
  FA_X1 u5_mult_82_S2_32_11 ( .A(u5_mult_82_ab_32__11_), .B(
        u5_mult_82_CARRYB_31__11_), .CI(u5_mult_82_SUMB_31__12_), .CO(
        u5_mult_82_CARRYB_32__11_), .S(u5_mult_82_SUMB_32__11_) );
  FA_X1 u5_mult_82_S2_32_10 ( .A(u5_mult_82_ab_32__10_), .B(
        u5_mult_82_CARRYB_31__10_), .CI(u5_mult_82_SUMB_31__11_), .CO(
        u5_mult_82_CARRYB_32__10_), .S(u5_mult_82_SUMB_32__10_) );
  FA_X1 u5_mult_82_S2_32_9 ( .A(u5_mult_82_ab_32__9_), .B(
        u5_mult_82_CARRYB_31__9_), .CI(u5_mult_82_SUMB_31__10_), .CO(
        u5_mult_82_CARRYB_32__9_), .S(u5_mult_82_SUMB_32__9_) );
  FA_X1 u5_mult_82_S2_32_8 ( .A(u5_mult_82_ab_32__8_), .B(
        u5_mult_82_CARRYB_31__8_), .CI(u5_mult_82_SUMB_31__9_), .CO(
        u5_mult_82_CARRYB_32__8_), .S(u5_mult_82_SUMB_32__8_) );
  FA_X1 u5_mult_82_S2_32_7 ( .A(u5_mult_82_ab_32__7_), .B(
        u5_mult_82_CARRYB_31__7_), .CI(u5_mult_82_SUMB_31__8_), .CO(
        u5_mult_82_CARRYB_32__7_), .S(u5_mult_82_SUMB_32__7_) );
  FA_X1 u5_mult_82_S2_32_6 ( .A(u5_mult_82_ab_32__6_), .B(
        u5_mult_82_CARRYB_31__6_), .CI(u5_mult_82_SUMB_31__7_), .CO(
        u5_mult_82_CARRYB_32__6_), .S(u5_mult_82_SUMB_32__6_) );
  FA_X1 u5_mult_82_S2_32_5 ( .A(u5_mult_82_ab_32__5_), .B(
        u5_mult_82_CARRYB_31__5_), .CI(u5_mult_82_SUMB_31__6_), .CO(
        u5_mult_82_CARRYB_32__5_), .S(u5_mult_82_SUMB_32__5_) );
  FA_X1 u5_mult_82_S2_32_4 ( .A(u5_mult_82_ab_32__4_), .B(
        u5_mult_82_CARRYB_31__4_), .CI(u5_mult_82_SUMB_31__5_), .CO(
        u5_mult_82_CARRYB_32__4_), .S(u5_mult_82_SUMB_32__4_) );
  FA_X1 u5_mult_82_S2_32_3 ( .A(u5_mult_82_ab_32__3_), .B(
        u5_mult_82_CARRYB_31__3_), .CI(u5_mult_82_SUMB_31__4_), .CO(
        u5_mult_82_CARRYB_32__3_), .S(u5_mult_82_SUMB_32__3_) );
  FA_X1 u5_mult_82_S2_32_2 ( .A(u5_mult_82_ab_32__2_), .B(
        u5_mult_82_CARRYB_31__2_), .CI(u5_mult_82_SUMB_31__3_), .CO(
        u5_mult_82_CARRYB_32__2_), .S(u5_mult_82_SUMB_32__2_) );
  FA_X1 u5_mult_82_S2_32_1 ( .A(u5_mult_82_ab_32__1_), .B(
        u5_mult_82_CARRYB_31__1_), .CI(u5_mult_82_SUMB_31__2_), .CO(
        u5_mult_82_CARRYB_32__1_), .S(u5_mult_82_SUMB_32__1_) );
  FA_X1 u5_mult_82_S1_32_0 ( .A(u5_mult_82_ab_32__0_), .B(
        u5_mult_82_CARRYB_31__0_), .CI(u5_mult_82_SUMB_31__1_), .CO(
        u5_mult_82_CARRYB_32__0_), .S(u5_N32) );
  FA_X1 u5_mult_82_S3_33_51 ( .A(u5_mult_82_ab_33__51_), .B(
        u5_mult_82_CARRYB_32__51_), .CI(u5_mult_82_ab_32__52_), .CO(
        u5_mult_82_CARRYB_33__51_), .S(u5_mult_82_SUMB_33__51_) );
  FA_X1 u5_mult_82_S2_33_50 ( .A(u5_mult_82_ab_33__50_), .B(
        u5_mult_82_CARRYB_32__50_), .CI(u5_mult_82_SUMB_32__51_), .CO(
        u5_mult_82_CARRYB_33__50_), .S(u5_mult_82_SUMB_33__50_) );
  FA_X1 u5_mult_82_S2_33_49 ( .A(u5_mult_82_ab_33__49_), .B(
        u5_mult_82_CARRYB_32__49_), .CI(u5_mult_82_SUMB_32__50_), .CO(
        u5_mult_82_CARRYB_33__49_), .S(u5_mult_82_SUMB_33__49_) );
  FA_X1 u5_mult_82_S2_33_48 ( .A(u5_mult_82_ab_33__48_), .B(
        u5_mult_82_CARRYB_32__48_), .CI(u5_mult_82_SUMB_32__49_), .CO(
        u5_mult_82_CARRYB_33__48_), .S(u5_mult_82_SUMB_33__48_) );
  FA_X1 u5_mult_82_S2_33_47 ( .A(u5_mult_82_ab_33__47_), .B(
        u5_mult_82_CARRYB_32__47_), .CI(u5_mult_82_SUMB_32__48_), .CO(
        u5_mult_82_CARRYB_33__47_), .S(u5_mult_82_SUMB_33__47_) );
  FA_X1 u5_mult_82_S2_33_46 ( .A(u5_mult_82_ab_33__46_), .B(
        u5_mult_82_CARRYB_32__46_), .CI(u5_mult_82_SUMB_32__47_), .CO(
        u5_mult_82_CARRYB_33__46_), .S(u5_mult_82_SUMB_33__46_) );
  FA_X1 u5_mult_82_S2_33_45 ( .A(u5_mult_82_ab_33__45_), .B(
        u5_mult_82_CARRYB_32__45_), .CI(u5_mult_82_SUMB_32__46_), .CO(
        u5_mult_82_CARRYB_33__45_), .S(u5_mult_82_SUMB_33__45_) );
  FA_X1 u5_mult_82_S2_33_44 ( .A(u5_mult_82_ab_33__44_), .B(
        u5_mult_82_CARRYB_32__44_), .CI(u5_mult_82_SUMB_32__45_), .CO(
        u5_mult_82_CARRYB_33__44_), .S(u5_mult_82_SUMB_33__44_) );
  FA_X1 u5_mult_82_S2_33_43 ( .A(u5_mult_82_ab_33__43_), .B(
        u5_mult_82_CARRYB_32__43_), .CI(u5_mult_82_SUMB_32__44_), .CO(
        u5_mult_82_CARRYB_33__43_), .S(u5_mult_82_SUMB_33__43_) );
  FA_X1 u5_mult_82_S2_33_42 ( .A(u5_mult_82_ab_33__42_), .B(
        u5_mult_82_CARRYB_32__42_), .CI(u5_mult_82_SUMB_32__43_), .CO(
        u5_mult_82_CARRYB_33__42_), .S(u5_mult_82_SUMB_33__42_) );
  FA_X1 u5_mult_82_S2_33_41 ( .A(u5_mult_82_ab_33__41_), .B(
        u5_mult_82_CARRYB_32__41_), .CI(u5_mult_82_SUMB_32__42_), .CO(
        u5_mult_82_CARRYB_33__41_), .S(u5_mult_82_SUMB_33__41_) );
  FA_X1 u5_mult_82_S2_33_40 ( .A(u5_mult_82_ab_33__40_), .B(
        u5_mult_82_CARRYB_32__40_), .CI(u5_mult_82_SUMB_32__41_), .CO(
        u5_mult_82_CARRYB_33__40_), .S(u5_mult_82_SUMB_33__40_) );
  FA_X1 u5_mult_82_S2_33_39 ( .A(u5_mult_82_ab_33__39_), .B(
        u5_mult_82_CARRYB_32__39_), .CI(u5_mult_82_SUMB_32__40_), .CO(
        u5_mult_82_CARRYB_33__39_), .S(u5_mult_82_SUMB_33__39_) );
  FA_X1 u5_mult_82_S2_33_38 ( .A(u5_mult_82_ab_33__38_), .B(
        u5_mult_82_CARRYB_32__38_), .CI(u5_mult_82_SUMB_32__39_), .CO(
        u5_mult_82_CARRYB_33__38_), .S(u5_mult_82_SUMB_33__38_) );
  FA_X1 u5_mult_82_S2_33_37 ( .A(u5_mult_82_ab_33__37_), .B(
        u5_mult_82_CARRYB_32__37_), .CI(u5_mult_82_SUMB_32__38_), .CO(
        u5_mult_82_CARRYB_33__37_), .S(u5_mult_82_SUMB_33__37_) );
  FA_X1 u5_mult_82_S2_33_36 ( .A(u5_mult_82_ab_33__36_), .B(
        u5_mult_82_CARRYB_32__36_), .CI(u5_mult_82_SUMB_32__37_), .CO(
        u5_mult_82_CARRYB_33__36_), .S(u5_mult_82_SUMB_33__36_) );
  FA_X1 u5_mult_82_S2_33_35 ( .A(u5_mult_82_ab_33__35_), .B(
        u5_mult_82_CARRYB_32__35_), .CI(u5_mult_82_SUMB_32__36_), .CO(
        u5_mult_82_CARRYB_33__35_), .S(u5_mult_82_SUMB_33__35_) );
  FA_X1 u5_mult_82_S2_33_34 ( .A(u5_mult_82_ab_33__34_), .B(
        u5_mult_82_CARRYB_32__34_), .CI(u5_mult_82_SUMB_32__35_), .CO(
        u5_mult_82_CARRYB_33__34_), .S(u5_mult_82_SUMB_33__34_) );
  FA_X1 u5_mult_82_S2_33_33 ( .A(u5_mult_82_ab_33__33_), .B(
        u5_mult_82_CARRYB_32__33_), .CI(u5_mult_82_SUMB_32__34_), .CO(
        u5_mult_82_CARRYB_33__33_), .S(u5_mult_82_SUMB_33__33_) );
  FA_X1 u5_mult_82_S2_33_32 ( .A(u5_mult_82_ab_33__32_), .B(
        u5_mult_82_CARRYB_32__32_), .CI(u5_mult_82_SUMB_32__33_), .CO(
        u5_mult_82_CARRYB_33__32_), .S(u5_mult_82_SUMB_33__32_) );
  FA_X1 u5_mult_82_S2_33_31 ( .A(u5_mult_82_ab_33__31_), .B(
        u5_mult_82_CARRYB_32__31_), .CI(u5_mult_82_SUMB_32__32_), .CO(
        u5_mult_82_CARRYB_33__31_), .S(u5_mult_82_SUMB_33__31_) );
  FA_X1 u5_mult_82_S2_33_30 ( .A(u5_mult_82_ab_33__30_), .B(
        u5_mult_82_CARRYB_32__30_), .CI(u5_mult_82_SUMB_32__31_), .CO(
        u5_mult_82_CARRYB_33__30_), .S(u5_mult_82_SUMB_33__30_) );
  FA_X1 u5_mult_82_S2_33_29 ( .A(u5_mult_82_ab_33__29_), .B(
        u5_mult_82_CARRYB_32__29_), .CI(u5_mult_82_SUMB_32__30_), .CO(
        u5_mult_82_CARRYB_33__29_), .S(u5_mult_82_SUMB_33__29_) );
  FA_X1 u5_mult_82_S2_33_28 ( .A(u5_mult_82_ab_33__28_), .B(
        u5_mult_82_CARRYB_32__28_), .CI(u5_mult_82_SUMB_32__29_), .CO(
        u5_mult_82_CARRYB_33__28_), .S(u5_mult_82_SUMB_33__28_) );
  FA_X1 u5_mult_82_S2_33_27 ( .A(u5_mult_82_ab_33__27_), .B(
        u5_mult_82_CARRYB_32__27_), .CI(u5_mult_82_SUMB_32__28_), .CO(
        u5_mult_82_CARRYB_33__27_), .S(u5_mult_82_SUMB_33__27_) );
  FA_X1 u5_mult_82_S2_33_26 ( .A(u5_mult_82_ab_33__26_), .B(
        u5_mult_82_CARRYB_32__26_), .CI(u5_mult_82_SUMB_32__27_), .CO(
        u5_mult_82_CARRYB_33__26_), .S(u5_mult_82_SUMB_33__26_) );
  FA_X1 u5_mult_82_S2_33_25 ( .A(u5_mult_82_ab_33__25_), .B(
        u5_mult_82_CARRYB_32__25_), .CI(u5_mult_82_SUMB_32__26_), .CO(
        u5_mult_82_CARRYB_33__25_), .S(u5_mult_82_SUMB_33__25_) );
  FA_X1 u5_mult_82_S2_33_24 ( .A(u5_mult_82_ab_33__24_), .B(
        u5_mult_82_CARRYB_32__24_), .CI(u5_mult_82_SUMB_32__25_), .CO(
        u5_mult_82_CARRYB_33__24_), .S(u5_mult_82_SUMB_33__24_) );
  FA_X1 u5_mult_82_S2_33_23 ( .A(u5_mult_82_ab_33__23_), .B(
        u5_mult_82_CARRYB_32__23_), .CI(u5_mult_82_SUMB_32__24_), .CO(
        u5_mult_82_CARRYB_33__23_), .S(u5_mult_82_SUMB_33__23_) );
  FA_X1 u5_mult_82_S2_33_22 ( .A(u5_mult_82_ab_33__22_), .B(
        u5_mult_82_CARRYB_32__22_), .CI(u5_mult_82_SUMB_32__23_), .CO(
        u5_mult_82_CARRYB_33__22_), .S(u5_mult_82_SUMB_33__22_) );
  FA_X1 u5_mult_82_S2_33_21 ( .A(u5_mult_82_ab_33__21_), .B(
        u5_mult_82_CARRYB_32__21_), .CI(u5_mult_82_SUMB_32__22_), .CO(
        u5_mult_82_CARRYB_33__21_), .S(u5_mult_82_SUMB_33__21_) );
  FA_X1 u5_mult_82_S2_33_20 ( .A(u5_mult_82_ab_33__20_), .B(
        u5_mult_82_CARRYB_32__20_), .CI(u5_mult_82_SUMB_32__21_), .CO(
        u5_mult_82_CARRYB_33__20_), .S(u5_mult_82_SUMB_33__20_) );
  FA_X1 u5_mult_82_S2_33_19 ( .A(u5_mult_82_ab_33__19_), .B(
        u5_mult_82_CARRYB_32__19_), .CI(u5_mult_82_SUMB_32__20_), .CO(
        u5_mult_82_CARRYB_33__19_), .S(u5_mult_82_SUMB_33__19_) );
  FA_X1 u5_mult_82_S2_33_18 ( .A(u5_mult_82_ab_33__18_), .B(
        u5_mult_82_CARRYB_32__18_), .CI(u5_mult_82_SUMB_32__19_), .CO(
        u5_mult_82_CARRYB_33__18_), .S(u5_mult_82_SUMB_33__18_) );
  FA_X1 u5_mult_82_S2_33_17 ( .A(u5_mult_82_ab_33__17_), .B(
        u5_mult_82_CARRYB_32__17_), .CI(u5_mult_82_SUMB_32__18_), .CO(
        u5_mult_82_CARRYB_33__17_), .S(u5_mult_82_SUMB_33__17_) );
  FA_X1 u5_mult_82_S2_33_16 ( .A(u5_mult_82_ab_33__16_), .B(
        u5_mult_82_CARRYB_32__16_), .CI(u5_mult_82_SUMB_32__17_), .CO(
        u5_mult_82_CARRYB_33__16_), .S(u5_mult_82_SUMB_33__16_) );
  FA_X1 u5_mult_82_S2_33_15 ( .A(u5_mult_82_ab_33__15_), .B(
        u5_mult_82_CARRYB_32__15_), .CI(u5_mult_82_SUMB_32__16_), .CO(
        u5_mult_82_CARRYB_33__15_), .S(u5_mult_82_SUMB_33__15_) );
  FA_X1 u5_mult_82_S2_33_14 ( .A(u5_mult_82_ab_33__14_), .B(
        u5_mult_82_CARRYB_32__14_), .CI(u5_mult_82_SUMB_32__15_), .CO(
        u5_mult_82_CARRYB_33__14_), .S(u5_mult_82_SUMB_33__14_) );
  FA_X1 u5_mult_82_S2_33_13 ( .A(u5_mult_82_ab_33__13_), .B(
        u5_mult_82_CARRYB_32__13_), .CI(u5_mult_82_SUMB_32__14_), .CO(
        u5_mult_82_CARRYB_33__13_), .S(u5_mult_82_SUMB_33__13_) );
  FA_X1 u5_mult_82_S2_33_12 ( .A(u5_mult_82_ab_33__12_), .B(
        u5_mult_82_CARRYB_32__12_), .CI(u5_mult_82_SUMB_32__13_), .CO(
        u5_mult_82_CARRYB_33__12_), .S(u5_mult_82_SUMB_33__12_) );
  FA_X1 u5_mult_82_S2_33_11 ( .A(u5_mult_82_ab_33__11_), .B(
        u5_mult_82_CARRYB_32__11_), .CI(u5_mult_82_SUMB_32__12_), .CO(
        u5_mult_82_CARRYB_33__11_), .S(u5_mult_82_SUMB_33__11_) );
  FA_X1 u5_mult_82_S2_33_10 ( .A(u5_mult_82_ab_33__10_), .B(
        u5_mult_82_CARRYB_32__10_), .CI(u5_mult_82_SUMB_32__11_), .CO(
        u5_mult_82_CARRYB_33__10_), .S(u5_mult_82_SUMB_33__10_) );
  FA_X1 u5_mult_82_S2_33_9 ( .A(u5_mult_82_ab_33__9_), .B(
        u5_mult_82_CARRYB_32__9_), .CI(u5_mult_82_SUMB_32__10_), .CO(
        u5_mult_82_CARRYB_33__9_), .S(u5_mult_82_SUMB_33__9_) );
  FA_X1 u5_mult_82_S2_33_8 ( .A(u5_mult_82_ab_33__8_), .B(
        u5_mult_82_CARRYB_32__8_), .CI(u5_mult_82_SUMB_32__9_), .CO(
        u5_mult_82_CARRYB_33__8_), .S(u5_mult_82_SUMB_33__8_) );
  FA_X1 u5_mult_82_S2_33_7 ( .A(u5_mult_82_ab_33__7_), .B(
        u5_mult_82_CARRYB_32__7_), .CI(u5_mult_82_SUMB_32__8_), .CO(
        u5_mult_82_CARRYB_33__7_), .S(u5_mult_82_SUMB_33__7_) );
  FA_X1 u5_mult_82_S2_33_6 ( .A(u5_mult_82_ab_33__6_), .B(
        u5_mult_82_CARRYB_32__6_), .CI(u5_mult_82_SUMB_32__7_), .CO(
        u5_mult_82_CARRYB_33__6_), .S(u5_mult_82_SUMB_33__6_) );
  FA_X1 u5_mult_82_S2_33_5 ( .A(u5_mult_82_ab_33__5_), .B(
        u5_mult_82_CARRYB_32__5_), .CI(u5_mult_82_SUMB_32__6_), .CO(
        u5_mult_82_CARRYB_33__5_), .S(u5_mult_82_SUMB_33__5_) );
  FA_X1 u5_mult_82_S2_33_4 ( .A(u5_mult_82_ab_33__4_), .B(
        u5_mult_82_CARRYB_32__4_), .CI(u5_mult_82_SUMB_32__5_), .CO(
        u5_mult_82_CARRYB_33__4_), .S(u5_mult_82_SUMB_33__4_) );
  FA_X1 u5_mult_82_S2_33_3 ( .A(u5_mult_82_ab_33__3_), .B(
        u5_mult_82_CARRYB_32__3_), .CI(u5_mult_82_SUMB_32__4_), .CO(
        u5_mult_82_CARRYB_33__3_), .S(u5_mult_82_SUMB_33__3_) );
  FA_X1 u5_mult_82_S2_33_2 ( .A(u5_mult_82_ab_33__2_), .B(
        u5_mult_82_CARRYB_32__2_), .CI(u5_mult_82_SUMB_32__3_), .CO(
        u5_mult_82_CARRYB_33__2_), .S(u5_mult_82_SUMB_33__2_) );
  FA_X1 u5_mult_82_S2_33_1 ( .A(u5_mult_82_ab_33__1_), .B(
        u5_mult_82_CARRYB_32__1_), .CI(u5_mult_82_SUMB_32__2_), .CO(
        u5_mult_82_CARRYB_33__1_), .S(u5_mult_82_SUMB_33__1_) );
  FA_X1 u5_mult_82_S1_33_0 ( .A(u5_mult_82_ab_33__0_), .B(
        u5_mult_82_CARRYB_32__0_), .CI(u5_mult_82_SUMB_32__1_), .CO(
        u5_mult_82_CARRYB_33__0_), .S(u5_N33) );
  FA_X1 u5_mult_82_S3_34_51 ( .A(u5_mult_82_ab_34__51_), .B(
        u5_mult_82_CARRYB_33__51_), .CI(u5_mult_82_ab_33__52_), .CO(
        u5_mult_82_CARRYB_34__51_), .S(u5_mult_82_SUMB_34__51_) );
  FA_X1 u5_mult_82_S2_34_50 ( .A(u5_mult_82_ab_34__50_), .B(
        u5_mult_82_CARRYB_33__50_), .CI(u5_mult_82_SUMB_33__51_), .CO(
        u5_mult_82_CARRYB_34__50_), .S(u5_mult_82_SUMB_34__50_) );
  FA_X1 u5_mult_82_S2_34_49 ( .A(u5_mult_82_ab_34__49_), .B(
        u5_mult_82_CARRYB_33__49_), .CI(u5_mult_82_SUMB_33__50_), .CO(
        u5_mult_82_CARRYB_34__49_), .S(u5_mult_82_SUMB_34__49_) );
  FA_X1 u5_mult_82_S2_34_48 ( .A(u5_mult_82_ab_34__48_), .B(
        u5_mult_82_CARRYB_33__48_), .CI(u5_mult_82_SUMB_33__49_), .CO(
        u5_mult_82_CARRYB_34__48_), .S(u5_mult_82_SUMB_34__48_) );
  FA_X1 u5_mult_82_S2_34_47 ( .A(u5_mult_82_ab_34__47_), .B(
        u5_mult_82_CARRYB_33__47_), .CI(u5_mult_82_SUMB_33__48_), .CO(
        u5_mult_82_CARRYB_34__47_), .S(u5_mult_82_SUMB_34__47_) );
  FA_X1 u5_mult_82_S2_34_46 ( .A(u5_mult_82_ab_34__46_), .B(
        u5_mult_82_CARRYB_33__46_), .CI(u5_mult_82_SUMB_33__47_), .CO(
        u5_mult_82_CARRYB_34__46_), .S(u5_mult_82_SUMB_34__46_) );
  FA_X1 u5_mult_82_S2_34_45 ( .A(u5_mult_82_ab_34__45_), .B(
        u5_mult_82_CARRYB_33__45_), .CI(u5_mult_82_SUMB_33__46_), .CO(
        u5_mult_82_CARRYB_34__45_), .S(u5_mult_82_SUMB_34__45_) );
  FA_X1 u5_mult_82_S2_34_44 ( .A(u5_mult_82_ab_34__44_), .B(
        u5_mult_82_CARRYB_33__44_), .CI(u5_mult_82_SUMB_33__45_), .CO(
        u5_mult_82_CARRYB_34__44_), .S(u5_mult_82_SUMB_34__44_) );
  FA_X1 u5_mult_82_S2_34_43 ( .A(u5_mult_82_ab_34__43_), .B(
        u5_mult_82_CARRYB_33__43_), .CI(u5_mult_82_SUMB_33__44_), .CO(
        u5_mult_82_CARRYB_34__43_), .S(u5_mult_82_SUMB_34__43_) );
  FA_X1 u5_mult_82_S2_34_42 ( .A(u5_mult_82_ab_34__42_), .B(
        u5_mult_82_CARRYB_33__42_), .CI(u5_mult_82_SUMB_33__43_), .CO(
        u5_mult_82_CARRYB_34__42_), .S(u5_mult_82_SUMB_34__42_) );
  FA_X1 u5_mult_82_S2_34_41 ( .A(u5_mult_82_ab_34__41_), .B(
        u5_mult_82_CARRYB_33__41_), .CI(u5_mult_82_SUMB_33__42_), .CO(
        u5_mult_82_CARRYB_34__41_), .S(u5_mult_82_SUMB_34__41_) );
  FA_X1 u5_mult_82_S2_34_40 ( .A(u5_mult_82_ab_34__40_), .B(
        u5_mult_82_CARRYB_33__40_), .CI(u5_mult_82_SUMB_33__41_), .CO(
        u5_mult_82_CARRYB_34__40_), .S(u5_mult_82_SUMB_34__40_) );
  FA_X1 u5_mult_82_S2_34_39 ( .A(u5_mult_82_ab_34__39_), .B(
        u5_mult_82_CARRYB_33__39_), .CI(u5_mult_82_SUMB_33__40_), .CO(
        u5_mult_82_CARRYB_34__39_), .S(u5_mult_82_SUMB_34__39_) );
  FA_X1 u5_mult_82_S2_34_38 ( .A(u5_mult_82_ab_34__38_), .B(
        u5_mult_82_CARRYB_33__38_), .CI(u5_mult_82_SUMB_33__39_), .CO(
        u5_mult_82_CARRYB_34__38_), .S(u5_mult_82_SUMB_34__38_) );
  FA_X1 u5_mult_82_S2_34_37 ( .A(u5_mult_82_ab_34__37_), .B(
        u5_mult_82_CARRYB_33__37_), .CI(u5_mult_82_SUMB_33__38_), .CO(
        u5_mult_82_CARRYB_34__37_), .S(u5_mult_82_SUMB_34__37_) );
  FA_X1 u5_mult_82_S2_34_36 ( .A(u5_mult_82_ab_34__36_), .B(
        u5_mult_82_CARRYB_33__36_), .CI(u5_mult_82_SUMB_33__37_), .CO(
        u5_mult_82_CARRYB_34__36_), .S(u5_mult_82_SUMB_34__36_) );
  FA_X1 u5_mult_82_S2_34_35 ( .A(u5_mult_82_ab_34__35_), .B(
        u5_mult_82_CARRYB_33__35_), .CI(u5_mult_82_SUMB_33__36_), .CO(
        u5_mult_82_CARRYB_34__35_), .S(u5_mult_82_SUMB_34__35_) );
  FA_X1 u5_mult_82_S2_34_34 ( .A(u5_mult_82_ab_34__34_), .B(
        u5_mult_82_CARRYB_33__34_), .CI(u5_mult_82_SUMB_33__35_), .CO(
        u5_mult_82_CARRYB_34__34_), .S(u5_mult_82_SUMB_34__34_) );
  FA_X1 u5_mult_82_S2_34_33 ( .A(u5_mult_82_ab_34__33_), .B(
        u5_mult_82_CARRYB_33__33_), .CI(u5_mult_82_SUMB_33__34_), .CO(
        u5_mult_82_CARRYB_34__33_), .S(u5_mult_82_SUMB_34__33_) );
  FA_X1 u5_mult_82_S2_34_32 ( .A(u5_mult_82_ab_34__32_), .B(
        u5_mult_82_CARRYB_33__32_), .CI(u5_mult_82_SUMB_33__33_), .CO(
        u5_mult_82_CARRYB_34__32_), .S(u5_mult_82_SUMB_34__32_) );
  FA_X1 u5_mult_82_S2_34_31 ( .A(u5_mult_82_ab_34__31_), .B(
        u5_mult_82_CARRYB_33__31_), .CI(u5_mult_82_SUMB_33__32_), .CO(
        u5_mult_82_CARRYB_34__31_), .S(u5_mult_82_SUMB_34__31_) );
  FA_X1 u5_mult_82_S2_34_30 ( .A(u5_mult_82_ab_34__30_), .B(
        u5_mult_82_CARRYB_33__30_), .CI(u5_mult_82_SUMB_33__31_), .CO(
        u5_mult_82_CARRYB_34__30_), .S(u5_mult_82_SUMB_34__30_) );
  FA_X1 u5_mult_82_S2_34_29 ( .A(u5_mult_82_ab_34__29_), .B(
        u5_mult_82_CARRYB_33__29_), .CI(u5_mult_82_SUMB_33__30_), .CO(
        u5_mult_82_CARRYB_34__29_), .S(u5_mult_82_SUMB_34__29_) );
  FA_X1 u5_mult_82_S2_34_28 ( .A(u5_mult_82_ab_34__28_), .B(
        u5_mult_82_CARRYB_33__28_), .CI(u5_mult_82_SUMB_33__29_), .CO(
        u5_mult_82_CARRYB_34__28_), .S(u5_mult_82_SUMB_34__28_) );
  FA_X1 u5_mult_82_S2_34_27 ( .A(u5_mult_82_ab_34__27_), .B(
        u5_mult_82_CARRYB_33__27_), .CI(u5_mult_82_SUMB_33__28_), .CO(
        u5_mult_82_CARRYB_34__27_), .S(u5_mult_82_SUMB_34__27_) );
  FA_X1 u5_mult_82_S2_34_26 ( .A(u5_mult_82_ab_34__26_), .B(
        u5_mult_82_CARRYB_33__26_), .CI(u5_mult_82_SUMB_33__27_), .CO(
        u5_mult_82_CARRYB_34__26_), .S(u5_mult_82_SUMB_34__26_) );
  FA_X1 u5_mult_82_S2_34_25 ( .A(u5_mult_82_ab_34__25_), .B(
        u5_mult_82_CARRYB_33__25_), .CI(u5_mult_82_SUMB_33__26_), .CO(
        u5_mult_82_CARRYB_34__25_), .S(u5_mult_82_SUMB_34__25_) );
  FA_X1 u5_mult_82_S2_34_24 ( .A(u5_mult_82_ab_34__24_), .B(
        u5_mult_82_CARRYB_33__24_), .CI(u5_mult_82_SUMB_33__25_), .CO(
        u5_mult_82_CARRYB_34__24_), .S(u5_mult_82_SUMB_34__24_) );
  FA_X1 u5_mult_82_S2_34_23 ( .A(u5_mult_82_ab_34__23_), .B(
        u5_mult_82_CARRYB_33__23_), .CI(u5_mult_82_SUMB_33__24_), .CO(
        u5_mult_82_CARRYB_34__23_), .S(u5_mult_82_SUMB_34__23_) );
  FA_X1 u5_mult_82_S2_34_22 ( .A(u5_mult_82_ab_34__22_), .B(
        u5_mult_82_CARRYB_33__22_), .CI(u5_mult_82_SUMB_33__23_), .CO(
        u5_mult_82_CARRYB_34__22_), .S(u5_mult_82_SUMB_34__22_) );
  FA_X1 u5_mult_82_S2_34_21 ( .A(u5_mult_82_ab_34__21_), .B(
        u5_mult_82_CARRYB_33__21_), .CI(u5_mult_82_SUMB_33__22_), .CO(
        u5_mult_82_CARRYB_34__21_), .S(u5_mult_82_SUMB_34__21_) );
  FA_X1 u5_mult_82_S2_34_20 ( .A(u5_mult_82_ab_34__20_), .B(
        u5_mult_82_CARRYB_33__20_), .CI(u5_mult_82_SUMB_33__21_), .CO(
        u5_mult_82_CARRYB_34__20_), .S(u5_mult_82_SUMB_34__20_) );
  FA_X1 u5_mult_82_S2_34_19 ( .A(u5_mult_82_ab_34__19_), .B(
        u5_mult_82_CARRYB_33__19_), .CI(u5_mult_82_SUMB_33__20_), .CO(
        u5_mult_82_CARRYB_34__19_), .S(u5_mult_82_SUMB_34__19_) );
  FA_X1 u5_mult_82_S2_34_18 ( .A(u5_mult_82_ab_34__18_), .B(
        u5_mult_82_CARRYB_33__18_), .CI(u5_mult_82_SUMB_33__19_), .CO(
        u5_mult_82_CARRYB_34__18_), .S(u5_mult_82_SUMB_34__18_) );
  FA_X1 u5_mult_82_S2_34_17 ( .A(u5_mult_82_ab_34__17_), .B(
        u5_mult_82_CARRYB_33__17_), .CI(u5_mult_82_SUMB_33__18_), .CO(
        u5_mult_82_CARRYB_34__17_), .S(u5_mult_82_SUMB_34__17_) );
  FA_X1 u5_mult_82_S2_34_16 ( .A(u5_mult_82_ab_34__16_), .B(
        u5_mult_82_CARRYB_33__16_), .CI(u5_mult_82_SUMB_33__17_), .CO(
        u5_mult_82_CARRYB_34__16_), .S(u5_mult_82_SUMB_34__16_) );
  FA_X1 u5_mult_82_S2_34_15 ( .A(u5_mult_82_ab_34__15_), .B(
        u5_mult_82_CARRYB_33__15_), .CI(u5_mult_82_SUMB_33__16_), .CO(
        u5_mult_82_CARRYB_34__15_), .S(u5_mult_82_SUMB_34__15_) );
  FA_X1 u5_mult_82_S2_34_14 ( .A(u5_mult_82_ab_34__14_), .B(
        u5_mult_82_CARRYB_33__14_), .CI(u5_mult_82_SUMB_33__15_), .CO(
        u5_mult_82_CARRYB_34__14_), .S(u5_mult_82_SUMB_34__14_) );
  FA_X1 u5_mult_82_S2_34_13 ( .A(u5_mult_82_ab_34__13_), .B(
        u5_mult_82_CARRYB_33__13_), .CI(u5_mult_82_SUMB_33__14_), .CO(
        u5_mult_82_CARRYB_34__13_), .S(u5_mult_82_SUMB_34__13_) );
  FA_X1 u5_mult_82_S2_34_12 ( .A(u5_mult_82_ab_34__12_), .B(
        u5_mult_82_CARRYB_33__12_), .CI(u5_mult_82_SUMB_33__13_), .CO(
        u5_mult_82_CARRYB_34__12_), .S(u5_mult_82_SUMB_34__12_) );
  FA_X1 u5_mult_82_S2_34_11 ( .A(u5_mult_82_ab_34__11_), .B(
        u5_mult_82_CARRYB_33__11_), .CI(u5_mult_82_SUMB_33__12_), .CO(
        u5_mult_82_CARRYB_34__11_), .S(u5_mult_82_SUMB_34__11_) );
  FA_X1 u5_mult_82_S2_34_10 ( .A(u5_mult_82_ab_34__10_), .B(
        u5_mult_82_CARRYB_33__10_), .CI(u5_mult_82_SUMB_33__11_), .CO(
        u5_mult_82_CARRYB_34__10_), .S(u5_mult_82_SUMB_34__10_) );
  FA_X1 u5_mult_82_S2_34_9 ( .A(u5_mult_82_ab_34__9_), .B(
        u5_mult_82_CARRYB_33__9_), .CI(u5_mult_82_SUMB_33__10_), .CO(
        u5_mult_82_CARRYB_34__9_), .S(u5_mult_82_SUMB_34__9_) );
  FA_X1 u5_mult_82_S2_34_8 ( .A(u5_mult_82_ab_34__8_), .B(
        u5_mult_82_CARRYB_33__8_), .CI(u5_mult_82_SUMB_33__9_), .CO(
        u5_mult_82_CARRYB_34__8_), .S(u5_mult_82_SUMB_34__8_) );
  FA_X1 u5_mult_82_S2_34_7 ( .A(u5_mult_82_ab_34__7_), .B(
        u5_mult_82_CARRYB_33__7_), .CI(u5_mult_82_SUMB_33__8_), .CO(
        u5_mult_82_CARRYB_34__7_), .S(u5_mult_82_SUMB_34__7_) );
  FA_X1 u5_mult_82_S2_34_6 ( .A(u5_mult_82_ab_34__6_), .B(
        u5_mult_82_CARRYB_33__6_), .CI(u5_mult_82_SUMB_33__7_), .CO(
        u5_mult_82_CARRYB_34__6_), .S(u5_mult_82_SUMB_34__6_) );
  FA_X1 u5_mult_82_S2_34_5 ( .A(u5_mult_82_ab_34__5_), .B(
        u5_mult_82_CARRYB_33__5_), .CI(u5_mult_82_SUMB_33__6_), .CO(
        u5_mult_82_CARRYB_34__5_), .S(u5_mult_82_SUMB_34__5_) );
  FA_X1 u5_mult_82_S2_34_4 ( .A(u5_mult_82_ab_34__4_), .B(
        u5_mult_82_CARRYB_33__4_), .CI(u5_mult_82_SUMB_33__5_), .CO(
        u5_mult_82_CARRYB_34__4_), .S(u5_mult_82_SUMB_34__4_) );
  FA_X1 u5_mult_82_S2_34_3 ( .A(u5_mult_82_ab_34__3_), .B(
        u5_mult_82_CARRYB_33__3_), .CI(u5_mult_82_SUMB_33__4_), .CO(
        u5_mult_82_CARRYB_34__3_), .S(u5_mult_82_SUMB_34__3_) );
  FA_X1 u5_mult_82_S2_34_2 ( .A(u5_mult_82_ab_34__2_), .B(
        u5_mult_82_CARRYB_33__2_), .CI(u5_mult_82_SUMB_33__3_), .CO(
        u5_mult_82_CARRYB_34__2_), .S(u5_mult_82_SUMB_34__2_) );
  FA_X1 u5_mult_82_S2_34_1 ( .A(u5_mult_82_ab_34__1_), .B(
        u5_mult_82_CARRYB_33__1_), .CI(u5_mult_82_SUMB_33__2_), .CO(
        u5_mult_82_CARRYB_34__1_), .S(u5_mult_82_SUMB_34__1_) );
  FA_X1 u5_mult_82_S1_34_0 ( .A(u5_mult_82_ab_34__0_), .B(
        u5_mult_82_CARRYB_33__0_), .CI(u5_mult_82_SUMB_33__1_), .CO(
        u5_mult_82_CARRYB_34__0_), .S(u5_N34) );
  FA_X1 u5_mult_82_S3_35_51 ( .A(u5_mult_82_ab_35__51_), .B(
        u5_mult_82_CARRYB_34__51_), .CI(u5_mult_82_ab_34__52_), .CO(
        u5_mult_82_CARRYB_35__51_), .S(u5_mult_82_SUMB_35__51_) );
  FA_X1 u5_mult_82_S2_35_50 ( .A(u5_mult_82_ab_35__50_), .B(
        u5_mult_82_CARRYB_34__50_), .CI(u5_mult_82_SUMB_34__51_), .CO(
        u5_mult_82_CARRYB_35__50_), .S(u5_mult_82_SUMB_35__50_) );
  FA_X1 u5_mult_82_S2_35_49 ( .A(u5_mult_82_ab_35__49_), .B(
        u5_mult_82_CARRYB_34__49_), .CI(u5_mult_82_SUMB_34__50_), .CO(
        u5_mult_82_CARRYB_35__49_), .S(u5_mult_82_SUMB_35__49_) );
  FA_X1 u5_mult_82_S2_35_48 ( .A(u5_mult_82_ab_35__48_), .B(
        u5_mult_82_CARRYB_34__48_), .CI(u5_mult_82_SUMB_34__49_), .CO(
        u5_mult_82_CARRYB_35__48_), .S(u5_mult_82_SUMB_35__48_) );
  FA_X1 u5_mult_82_S2_35_47 ( .A(u5_mult_82_ab_35__47_), .B(
        u5_mult_82_CARRYB_34__47_), .CI(u5_mult_82_SUMB_34__48_), .CO(
        u5_mult_82_CARRYB_35__47_), .S(u5_mult_82_SUMB_35__47_) );
  FA_X1 u5_mult_82_S2_35_46 ( .A(u5_mult_82_ab_35__46_), .B(
        u5_mult_82_CARRYB_34__46_), .CI(u5_mult_82_SUMB_34__47_), .CO(
        u5_mult_82_CARRYB_35__46_), .S(u5_mult_82_SUMB_35__46_) );
  FA_X1 u5_mult_82_S2_35_45 ( .A(u5_mult_82_ab_35__45_), .B(
        u5_mult_82_CARRYB_34__45_), .CI(u5_mult_82_SUMB_34__46_), .CO(
        u5_mult_82_CARRYB_35__45_), .S(u5_mult_82_SUMB_35__45_) );
  FA_X1 u5_mult_82_S2_35_44 ( .A(u5_mult_82_ab_35__44_), .B(
        u5_mult_82_CARRYB_34__44_), .CI(u5_mult_82_SUMB_34__45_), .CO(
        u5_mult_82_CARRYB_35__44_), .S(u5_mult_82_SUMB_35__44_) );
  FA_X1 u5_mult_82_S2_35_43 ( .A(u5_mult_82_ab_35__43_), .B(
        u5_mult_82_CARRYB_34__43_), .CI(u5_mult_82_SUMB_34__44_), .CO(
        u5_mult_82_CARRYB_35__43_), .S(u5_mult_82_SUMB_35__43_) );
  FA_X1 u5_mult_82_S2_35_42 ( .A(u5_mult_82_ab_35__42_), .B(
        u5_mult_82_CARRYB_34__42_), .CI(u5_mult_82_SUMB_34__43_), .CO(
        u5_mult_82_CARRYB_35__42_), .S(u5_mult_82_SUMB_35__42_) );
  FA_X1 u5_mult_82_S2_35_41 ( .A(u5_mult_82_ab_35__41_), .B(
        u5_mult_82_CARRYB_34__41_), .CI(u5_mult_82_SUMB_34__42_), .CO(
        u5_mult_82_CARRYB_35__41_), .S(u5_mult_82_SUMB_35__41_) );
  FA_X1 u5_mult_82_S2_35_40 ( .A(u5_mult_82_ab_35__40_), .B(
        u5_mult_82_CARRYB_34__40_), .CI(u5_mult_82_SUMB_34__41_), .CO(
        u5_mult_82_CARRYB_35__40_), .S(u5_mult_82_SUMB_35__40_) );
  FA_X1 u5_mult_82_S2_35_39 ( .A(u5_mult_82_ab_35__39_), .B(
        u5_mult_82_CARRYB_34__39_), .CI(u5_mult_82_SUMB_34__40_), .CO(
        u5_mult_82_CARRYB_35__39_), .S(u5_mult_82_SUMB_35__39_) );
  FA_X1 u5_mult_82_S2_35_38 ( .A(u5_mult_82_ab_35__38_), .B(
        u5_mult_82_CARRYB_34__38_), .CI(u5_mult_82_SUMB_34__39_), .CO(
        u5_mult_82_CARRYB_35__38_), .S(u5_mult_82_SUMB_35__38_) );
  FA_X1 u5_mult_82_S2_35_37 ( .A(u5_mult_82_ab_35__37_), .B(
        u5_mult_82_CARRYB_34__37_), .CI(u5_mult_82_SUMB_34__38_), .CO(
        u5_mult_82_CARRYB_35__37_), .S(u5_mult_82_SUMB_35__37_) );
  FA_X1 u5_mult_82_S2_35_36 ( .A(u5_mult_82_ab_35__36_), .B(
        u5_mult_82_CARRYB_34__36_), .CI(u5_mult_82_SUMB_34__37_), .CO(
        u5_mult_82_CARRYB_35__36_), .S(u5_mult_82_SUMB_35__36_) );
  FA_X1 u5_mult_82_S2_35_35 ( .A(u5_mult_82_ab_35__35_), .B(
        u5_mult_82_CARRYB_34__35_), .CI(u5_mult_82_SUMB_34__36_), .CO(
        u5_mult_82_CARRYB_35__35_), .S(u5_mult_82_SUMB_35__35_) );
  FA_X1 u5_mult_82_S2_35_34 ( .A(u5_mult_82_ab_35__34_), .B(
        u5_mult_82_CARRYB_34__34_), .CI(u5_mult_82_SUMB_34__35_), .CO(
        u5_mult_82_CARRYB_35__34_), .S(u5_mult_82_SUMB_35__34_) );
  FA_X1 u5_mult_82_S2_35_33 ( .A(u5_mult_82_ab_35__33_), .B(
        u5_mult_82_CARRYB_34__33_), .CI(u5_mult_82_SUMB_34__34_), .CO(
        u5_mult_82_CARRYB_35__33_), .S(u5_mult_82_SUMB_35__33_) );
  FA_X1 u5_mult_82_S2_35_32 ( .A(u5_mult_82_ab_35__32_), .B(
        u5_mult_82_CARRYB_34__32_), .CI(u5_mult_82_SUMB_34__33_), .CO(
        u5_mult_82_CARRYB_35__32_), .S(u5_mult_82_SUMB_35__32_) );
  FA_X1 u5_mult_82_S2_35_31 ( .A(u5_mult_82_ab_35__31_), .B(
        u5_mult_82_CARRYB_34__31_), .CI(u5_mult_82_SUMB_34__32_), .CO(
        u5_mult_82_CARRYB_35__31_), .S(u5_mult_82_SUMB_35__31_) );
  FA_X1 u5_mult_82_S2_35_30 ( .A(u5_mult_82_ab_35__30_), .B(
        u5_mult_82_CARRYB_34__30_), .CI(u5_mult_82_SUMB_34__31_), .CO(
        u5_mult_82_CARRYB_35__30_), .S(u5_mult_82_SUMB_35__30_) );
  FA_X1 u5_mult_82_S2_35_29 ( .A(u5_mult_82_ab_35__29_), .B(
        u5_mult_82_CARRYB_34__29_), .CI(u5_mult_82_SUMB_34__30_), .CO(
        u5_mult_82_CARRYB_35__29_), .S(u5_mult_82_SUMB_35__29_) );
  FA_X1 u5_mult_82_S2_35_28 ( .A(u5_mult_82_ab_35__28_), .B(
        u5_mult_82_CARRYB_34__28_), .CI(u5_mult_82_SUMB_34__29_), .CO(
        u5_mult_82_CARRYB_35__28_), .S(u5_mult_82_SUMB_35__28_) );
  FA_X1 u5_mult_82_S2_35_27 ( .A(u5_mult_82_ab_35__27_), .B(
        u5_mult_82_CARRYB_34__27_), .CI(u5_mult_82_SUMB_34__28_), .CO(
        u5_mult_82_CARRYB_35__27_), .S(u5_mult_82_SUMB_35__27_) );
  FA_X1 u5_mult_82_S2_35_26 ( .A(u5_mult_82_ab_35__26_), .B(
        u5_mult_82_CARRYB_34__26_), .CI(u5_mult_82_SUMB_34__27_), .CO(
        u5_mult_82_CARRYB_35__26_), .S(u5_mult_82_SUMB_35__26_) );
  FA_X1 u5_mult_82_S2_35_25 ( .A(u5_mult_82_ab_35__25_), .B(
        u5_mult_82_CARRYB_34__25_), .CI(u5_mult_82_SUMB_34__26_), .CO(
        u5_mult_82_CARRYB_35__25_), .S(u5_mult_82_SUMB_35__25_) );
  FA_X1 u5_mult_82_S2_35_24 ( .A(u5_mult_82_ab_35__24_), .B(
        u5_mult_82_CARRYB_34__24_), .CI(u5_mult_82_SUMB_34__25_), .CO(
        u5_mult_82_CARRYB_35__24_), .S(u5_mult_82_SUMB_35__24_) );
  FA_X1 u5_mult_82_S2_35_23 ( .A(u5_mult_82_ab_35__23_), .B(
        u5_mult_82_CARRYB_34__23_), .CI(u5_mult_82_SUMB_34__24_), .CO(
        u5_mult_82_CARRYB_35__23_), .S(u5_mult_82_SUMB_35__23_) );
  FA_X1 u5_mult_82_S2_35_22 ( .A(u5_mult_82_ab_35__22_), .B(
        u5_mult_82_CARRYB_34__22_), .CI(u5_mult_82_SUMB_34__23_), .CO(
        u5_mult_82_CARRYB_35__22_), .S(u5_mult_82_SUMB_35__22_) );
  FA_X1 u5_mult_82_S2_35_21 ( .A(u5_mult_82_ab_35__21_), .B(
        u5_mult_82_CARRYB_34__21_), .CI(u5_mult_82_SUMB_34__22_), .CO(
        u5_mult_82_CARRYB_35__21_), .S(u5_mult_82_SUMB_35__21_) );
  FA_X1 u5_mult_82_S2_35_20 ( .A(u5_mult_82_ab_35__20_), .B(
        u5_mult_82_CARRYB_34__20_), .CI(u5_mult_82_SUMB_34__21_), .CO(
        u5_mult_82_CARRYB_35__20_), .S(u5_mult_82_SUMB_35__20_) );
  FA_X1 u5_mult_82_S2_35_19 ( .A(u5_mult_82_ab_35__19_), .B(
        u5_mult_82_CARRYB_34__19_), .CI(u5_mult_82_SUMB_34__20_), .CO(
        u5_mult_82_CARRYB_35__19_), .S(u5_mult_82_SUMB_35__19_) );
  FA_X1 u5_mult_82_S2_35_18 ( .A(u5_mult_82_ab_35__18_), .B(
        u5_mult_82_CARRYB_34__18_), .CI(u5_mult_82_SUMB_34__19_), .CO(
        u5_mult_82_CARRYB_35__18_), .S(u5_mult_82_SUMB_35__18_) );
  FA_X1 u5_mult_82_S2_35_17 ( .A(u5_mult_82_ab_35__17_), .B(
        u5_mult_82_CARRYB_34__17_), .CI(u5_mult_82_SUMB_34__18_), .CO(
        u5_mult_82_CARRYB_35__17_), .S(u5_mult_82_SUMB_35__17_) );
  FA_X1 u5_mult_82_S2_35_16 ( .A(u5_mult_82_ab_35__16_), .B(
        u5_mult_82_CARRYB_34__16_), .CI(u5_mult_82_SUMB_34__17_), .CO(
        u5_mult_82_CARRYB_35__16_), .S(u5_mult_82_SUMB_35__16_) );
  FA_X1 u5_mult_82_S2_35_15 ( .A(u5_mult_82_ab_35__15_), .B(
        u5_mult_82_CARRYB_34__15_), .CI(u5_mult_82_SUMB_34__16_), .CO(
        u5_mult_82_CARRYB_35__15_), .S(u5_mult_82_SUMB_35__15_) );
  FA_X1 u5_mult_82_S2_35_14 ( .A(u5_mult_82_ab_35__14_), .B(
        u5_mult_82_CARRYB_34__14_), .CI(u5_mult_82_SUMB_34__15_), .CO(
        u5_mult_82_CARRYB_35__14_), .S(u5_mult_82_SUMB_35__14_) );
  FA_X1 u5_mult_82_S2_35_13 ( .A(u5_mult_82_ab_35__13_), .B(
        u5_mult_82_CARRYB_34__13_), .CI(u5_mult_82_SUMB_34__14_), .CO(
        u5_mult_82_CARRYB_35__13_), .S(u5_mult_82_SUMB_35__13_) );
  FA_X1 u5_mult_82_S2_35_12 ( .A(u5_mult_82_ab_35__12_), .B(
        u5_mult_82_CARRYB_34__12_), .CI(u5_mult_82_SUMB_34__13_), .CO(
        u5_mult_82_CARRYB_35__12_), .S(u5_mult_82_SUMB_35__12_) );
  FA_X1 u5_mult_82_S2_35_11 ( .A(u5_mult_82_ab_35__11_), .B(
        u5_mult_82_CARRYB_34__11_), .CI(u5_mult_82_SUMB_34__12_), .CO(
        u5_mult_82_CARRYB_35__11_), .S(u5_mult_82_SUMB_35__11_) );
  FA_X1 u5_mult_82_S2_35_10 ( .A(u5_mult_82_ab_35__10_), .B(
        u5_mult_82_CARRYB_34__10_), .CI(u5_mult_82_SUMB_34__11_), .CO(
        u5_mult_82_CARRYB_35__10_), .S(u5_mult_82_SUMB_35__10_) );
  FA_X1 u5_mult_82_S2_35_9 ( .A(u5_mult_82_ab_35__9_), .B(
        u5_mult_82_CARRYB_34__9_), .CI(u5_mult_82_SUMB_34__10_), .CO(
        u5_mult_82_CARRYB_35__9_), .S(u5_mult_82_SUMB_35__9_) );
  FA_X1 u5_mult_82_S2_35_8 ( .A(u5_mult_82_ab_35__8_), .B(
        u5_mult_82_CARRYB_34__8_), .CI(u5_mult_82_SUMB_34__9_), .CO(
        u5_mult_82_CARRYB_35__8_), .S(u5_mult_82_SUMB_35__8_) );
  FA_X1 u5_mult_82_S2_35_7 ( .A(u5_mult_82_ab_35__7_), .B(
        u5_mult_82_CARRYB_34__7_), .CI(u5_mult_82_SUMB_34__8_), .CO(
        u5_mult_82_CARRYB_35__7_), .S(u5_mult_82_SUMB_35__7_) );
  FA_X1 u5_mult_82_S2_35_6 ( .A(u5_mult_82_ab_35__6_), .B(
        u5_mult_82_CARRYB_34__6_), .CI(u5_mult_82_SUMB_34__7_), .CO(
        u5_mult_82_CARRYB_35__6_), .S(u5_mult_82_SUMB_35__6_) );
  FA_X1 u5_mult_82_S2_35_5 ( .A(u5_mult_82_ab_35__5_), .B(
        u5_mult_82_CARRYB_34__5_), .CI(u5_mult_82_SUMB_34__6_), .CO(
        u5_mult_82_CARRYB_35__5_), .S(u5_mult_82_SUMB_35__5_) );
  FA_X1 u5_mult_82_S2_35_4 ( .A(u5_mult_82_ab_35__4_), .B(
        u5_mult_82_CARRYB_34__4_), .CI(u5_mult_82_SUMB_34__5_), .CO(
        u5_mult_82_CARRYB_35__4_), .S(u5_mult_82_SUMB_35__4_) );
  FA_X1 u5_mult_82_S2_35_3 ( .A(u5_mult_82_ab_35__3_), .B(
        u5_mult_82_CARRYB_34__3_), .CI(u5_mult_82_SUMB_34__4_), .CO(
        u5_mult_82_CARRYB_35__3_), .S(u5_mult_82_SUMB_35__3_) );
  FA_X1 u5_mult_82_S2_35_2 ( .A(u5_mult_82_ab_35__2_), .B(
        u5_mult_82_CARRYB_34__2_), .CI(u5_mult_82_SUMB_34__3_), .CO(
        u5_mult_82_CARRYB_35__2_), .S(u5_mult_82_SUMB_35__2_) );
  FA_X1 u5_mult_82_S2_35_1 ( .A(u5_mult_82_ab_35__1_), .B(
        u5_mult_82_CARRYB_34__1_), .CI(u5_mult_82_SUMB_34__2_), .CO(
        u5_mult_82_CARRYB_35__1_), .S(u5_mult_82_SUMB_35__1_) );
  FA_X1 u5_mult_82_S1_35_0 ( .A(u5_mult_82_ab_35__0_), .B(
        u5_mult_82_CARRYB_34__0_), .CI(u5_mult_82_SUMB_34__1_), .CO(
        u5_mult_82_CARRYB_35__0_), .S(u5_N35) );
  FA_X1 u5_mult_82_S3_36_51 ( .A(u5_mult_82_ab_36__51_), .B(
        u5_mult_82_CARRYB_35__51_), .CI(u5_mult_82_ab_35__52_), .CO(
        u5_mult_82_CARRYB_36__51_), .S(u5_mult_82_SUMB_36__51_) );
  FA_X1 u5_mult_82_S2_36_50 ( .A(u5_mult_82_ab_36__50_), .B(
        u5_mult_82_CARRYB_35__50_), .CI(u5_mult_82_SUMB_35__51_), .CO(
        u5_mult_82_CARRYB_36__50_), .S(u5_mult_82_SUMB_36__50_) );
  FA_X1 u5_mult_82_S2_36_49 ( .A(u5_mult_82_ab_36__49_), .B(
        u5_mult_82_CARRYB_35__49_), .CI(u5_mult_82_SUMB_35__50_), .CO(
        u5_mult_82_CARRYB_36__49_), .S(u5_mult_82_SUMB_36__49_) );
  FA_X1 u5_mult_82_S2_36_48 ( .A(u5_mult_82_ab_36__48_), .B(
        u5_mult_82_CARRYB_35__48_), .CI(u5_mult_82_SUMB_35__49_), .CO(
        u5_mult_82_CARRYB_36__48_), .S(u5_mult_82_SUMB_36__48_) );
  FA_X1 u5_mult_82_S2_36_47 ( .A(u5_mult_82_ab_36__47_), .B(
        u5_mult_82_CARRYB_35__47_), .CI(u5_mult_82_SUMB_35__48_), .CO(
        u5_mult_82_CARRYB_36__47_), .S(u5_mult_82_SUMB_36__47_) );
  FA_X1 u5_mult_82_S2_36_46 ( .A(u5_mult_82_ab_36__46_), .B(
        u5_mult_82_CARRYB_35__46_), .CI(u5_mult_82_SUMB_35__47_), .CO(
        u5_mult_82_CARRYB_36__46_), .S(u5_mult_82_SUMB_36__46_) );
  FA_X1 u5_mult_82_S2_36_45 ( .A(u5_mult_82_ab_36__45_), .B(
        u5_mult_82_CARRYB_35__45_), .CI(u5_mult_82_SUMB_35__46_), .CO(
        u5_mult_82_CARRYB_36__45_), .S(u5_mult_82_SUMB_36__45_) );
  FA_X1 u5_mult_82_S2_36_44 ( .A(u5_mult_82_ab_36__44_), .B(
        u5_mult_82_CARRYB_35__44_), .CI(u5_mult_82_SUMB_35__45_), .CO(
        u5_mult_82_CARRYB_36__44_), .S(u5_mult_82_SUMB_36__44_) );
  FA_X1 u5_mult_82_S2_36_43 ( .A(u5_mult_82_ab_36__43_), .B(
        u5_mult_82_CARRYB_35__43_), .CI(u5_mult_82_SUMB_35__44_), .CO(
        u5_mult_82_CARRYB_36__43_), .S(u5_mult_82_SUMB_36__43_) );
  FA_X1 u5_mult_82_S2_36_42 ( .A(u5_mult_82_ab_36__42_), .B(
        u5_mult_82_CARRYB_35__42_), .CI(u5_mult_82_SUMB_35__43_), .CO(
        u5_mult_82_CARRYB_36__42_), .S(u5_mult_82_SUMB_36__42_) );
  FA_X1 u5_mult_82_S2_36_41 ( .A(u5_mult_82_ab_36__41_), .B(
        u5_mult_82_CARRYB_35__41_), .CI(u5_mult_82_SUMB_35__42_), .CO(
        u5_mult_82_CARRYB_36__41_), .S(u5_mult_82_SUMB_36__41_) );
  FA_X1 u5_mult_82_S2_36_40 ( .A(u5_mult_82_ab_36__40_), .B(
        u5_mult_82_CARRYB_35__40_), .CI(u5_mult_82_SUMB_35__41_), .CO(
        u5_mult_82_CARRYB_36__40_), .S(u5_mult_82_SUMB_36__40_) );
  FA_X1 u5_mult_82_S2_36_39 ( .A(u5_mult_82_ab_36__39_), .B(
        u5_mult_82_CARRYB_35__39_), .CI(u5_mult_82_SUMB_35__40_), .CO(
        u5_mult_82_CARRYB_36__39_), .S(u5_mult_82_SUMB_36__39_) );
  FA_X1 u5_mult_82_S2_36_38 ( .A(u5_mult_82_ab_36__38_), .B(
        u5_mult_82_CARRYB_35__38_), .CI(u5_mult_82_SUMB_35__39_), .CO(
        u5_mult_82_CARRYB_36__38_), .S(u5_mult_82_SUMB_36__38_) );
  FA_X1 u5_mult_82_S2_36_37 ( .A(u5_mult_82_ab_36__37_), .B(
        u5_mult_82_CARRYB_35__37_), .CI(u5_mult_82_SUMB_35__38_), .CO(
        u5_mult_82_CARRYB_36__37_), .S(u5_mult_82_SUMB_36__37_) );
  FA_X1 u5_mult_82_S2_36_36 ( .A(u5_mult_82_ab_36__36_), .B(
        u5_mult_82_CARRYB_35__36_), .CI(u5_mult_82_SUMB_35__37_), .CO(
        u5_mult_82_CARRYB_36__36_), .S(u5_mult_82_SUMB_36__36_) );
  FA_X1 u5_mult_82_S2_36_35 ( .A(u5_mult_82_ab_36__35_), .B(
        u5_mult_82_CARRYB_35__35_), .CI(u5_mult_82_SUMB_35__36_), .CO(
        u5_mult_82_CARRYB_36__35_), .S(u5_mult_82_SUMB_36__35_) );
  FA_X1 u5_mult_82_S2_36_34 ( .A(u5_mult_82_ab_36__34_), .B(
        u5_mult_82_CARRYB_35__34_), .CI(u5_mult_82_SUMB_35__35_), .CO(
        u5_mult_82_CARRYB_36__34_), .S(u5_mult_82_SUMB_36__34_) );
  FA_X1 u5_mult_82_S2_36_33 ( .A(u5_mult_82_ab_36__33_), .B(
        u5_mult_82_CARRYB_35__33_), .CI(u5_mult_82_SUMB_35__34_), .CO(
        u5_mult_82_CARRYB_36__33_), .S(u5_mult_82_SUMB_36__33_) );
  FA_X1 u5_mult_82_S2_36_32 ( .A(u5_mult_82_ab_36__32_), .B(
        u5_mult_82_CARRYB_35__32_), .CI(u5_mult_82_SUMB_35__33_), .CO(
        u5_mult_82_CARRYB_36__32_), .S(u5_mult_82_SUMB_36__32_) );
  FA_X1 u5_mult_82_S2_36_31 ( .A(u5_mult_82_ab_36__31_), .B(
        u5_mult_82_CARRYB_35__31_), .CI(u5_mult_82_SUMB_35__32_), .CO(
        u5_mult_82_CARRYB_36__31_), .S(u5_mult_82_SUMB_36__31_) );
  FA_X1 u5_mult_82_S2_36_30 ( .A(u5_mult_82_ab_36__30_), .B(
        u5_mult_82_CARRYB_35__30_), .CI(u5_mult_82_SUMB_35__31_), .CO(
        u5_mult_82_CARRYB_36__30_), .S(u5_mult_82_SUMB_36__30_) );
  FA_X1 u5_mult_82_S2_36_29 ( .A(u5_mult_82_ab_36__29_), .B(
        u5_mult_82_CARRYB_35__29_), .CI(u5_mult_82_SUMB_35__30_), .CO(
        u5_mult_82_CARRYB_36__29_), .S(u5_mult_82_SUMB_36__29_) );
  FA_X1 u5_mult_82_S2_36_28 ( .A(u5_mult_82_ab_36__28_), .B(
        u5_mult_82_CARRYB_35__28_), .CI(u5_mult_82_SUMB_35__29_), .CO(
        u5_mult_82_CARRYB_36__28_), .S(u5_mult_82_SUMB_36__28_) );
  FA_X1 u5_mult_82_S2_36_27 ( .A(u5_mult_82_ab_36__27_), .B(
        u5_mult_82_CARRYB_35__27_), .CI(u5_mult_82_SUMB_35__28_), .CO(
        u5_mult_82_CARRYB_36__27_), .S(u5_mult_82_SUMB_36__27_) );
  FA_X1 u5_mult_82_S2_36_26 ( .A(u5_mult_82_ab_36__26_), .B(
        u5_mult_82_CARRYB_35__26_), .CI(u5_mult_82_SUMB_35__27_), .CO(
        u5_mult_82_CARRYB_36__26_), .S(u5_mult_82_SUMB_36__26_) );
  FA_X1 u5_mult_82_S2_36_25 ( .A(u5_mult_82_ab_36__25_), .B(
        u5_mult_82_CARRYB_35__25_), .CI(u5_mult_82_SUMB_35__26_), .CO(
        u5_mult_82_CARRYB_36__25_), .S(u5_mult_82_SUMB_36__25_) );
  FA_X1 u5_mult_82_S2_36_24 ( .A(u5_mult_82_ab_36__24_), .B(
        u5_mult_82_CARRYB_35__24_), .CI(u5_mult_82_SUMB_35__25_), .CO(
        u5_mult_82_CARRYB_36__24_), .S(u5_mult_82_SUMB_36__24_) );
  FA_X1 u5_mult_82_S2_36_23 ( .A(u5_mult_82_ab_36__23_), .B(
        u5_mult_82_CARRYB_35__23_), .CI(u5_mult_82_SUMB_35__24_), .CO(
        u5_mult_82_CARRYB_36__23_), .S(u5_mult_82_SUMB_36__23_) );
  FA_X1 u5_mult_82_S2_36_22 ( .A(u5_mult_82_ab_36__22_), .B(
        u5_mult_82_CARRYB_35__22_), .CI(u5_mult_82_SUMB_35__23_), .CO(
        u5_mult_82_CARRYB_36__22_), .S(u5_mult_82_SUMB_36__22_) );
  FA_X1 u5_mult_82_S2_36_21 ( .A(u5_mult_82_ab_36__21_), .B(
        u5_mult_82_CARRYB_35__21_), .CI(u5_mult_82_SUMB_35__22_), .CO(
        u5_mult_82_CARRYB_36__21_), .S(u5_mult_82_SUMB_36__21_) );
  FA_X1 u5_mult_82_S2_36_20 ( .A(u5_mult_82_ab_36__20_), .B(
        u5_mult_82_CARRYB_35__20_), .CI(u5_mult_82_SUMB_35__21_), .CO(
        u5_mult_82_CARRYB_36__20_), .S(u5_mult_82_SUMB_36__20_) );
  FA_X1 u5_mult_82_S2_36_19 ( .A(u5_mult_82_ab_36__19_), .B(
        u5_mult_82_CARRYB_35__19_), .CI(u5_mult_82_SUMB_35__20_), .CO(
        u5_mult_82_CARRYB_36__19_), .S(u5_mult_82_SUMB_36__19_) );
  FA_X1 u5_mult_82_S2_36_18 ( .A(u5_mult_82_ab_36__18_), .B(
        u5_mult_82_CARRYB_35__18_), .CI(u5_mult_82_SUMB_35__19_), .CO(
        u5_mult_82_CARRYB_36__18_), .S(u5_mult_82_SUMB_36__18_) );
  FA_X1 u5_mult_82_S2_36_17 ( .A(u5_mult_82_ab_36__17_), .B(
        u5_mult_82_CARRYB_35__17_), .CI(u5_mult_82_SUMB_35__18_), .CO(
        u5_mult_82_CARRYB_36__17_), .S(u5_mult_82_SUMB_36__17_) );
  FA_X1 u5_mult_82_S2_36_16 ( .A(u5_mult_82_ab_36__16_), .B(
        u5_mult_82_CARRYB_35__16_), .CI(u5_mult_82_SUMB_35__17_), .CO(
        u5_mult_82_CARRYB_36__16_), .S(u5_mult_82_SUMB_36__16_) );
  FA_X1 u5_mult_82_S2_36_15 ( .A(u5_mult_82_ab_36__15_), .B(
        u5_mult_82_CARRYB_35__15_), .CI(u5_mult_82_SUMB_35__16_), .CO(
        u5_mult_82_CARRYB_36__15_), .S(u5_mult_82_SUMB_36__15_) );
  FA_X1 u5_mult_82_S2_36_14 ( .A(u5_mult_82_ab_36__14_), .B(
        u5_mult_82_CARRYB_35__14_), .CI(u5_mult_82_SUMB_35__15_), .CO(
        u5_mult_82_CARRYB_36__14_), .S(u5_mult_82_SUMB_36__14_) );
  FA_X1 u5_mult_82_S2_36_13 ( .A(u5_mult_82_ab_36__13_), .B(
        u5_mult_82_CARRYB_35__13_), .CI(u5_mult_82_SUMB_35__14_), .CO(
        u5_mult_82_CARRYB_36__13_), .S(u5_mult_82_SUMB_36__13_) );
  FA_X1 u5_mult_82_S2_36_12 ( .A(u5_mult_82_ab_36__12_), .B(
        u5_mult_82_CARRYB_35__12_), .CI(u5_mult_82_SUMB_35__13_), .CO(
        u5_mult_82_CARRYB_36__12_), .S(u5_mult_82_SUMB_36__12_) );
  FA_X1 u5_mult_82_S2_36_11 ( .A(u5_mult_82_ab_36__11_), .B(
        u5_mult_82_CARRYB_35__11_), .CI(u5_mult_82_SUMB_35__12_), .CO(
        u5_mult_82_CARRYB_36__11_), .S(u5_mult_82_SUMB_36__11_) );
  FA_X1 u5_mult_82_S2_36_10 ( .A(u5_mult_82_ab_36__10_), .B(
        u5_mult_82_CARRYB_35__10_), .CI(u5_mult_82_SUMB_35__11_), .CO(
        u5_mult_82_CARRYB_36__10_), .S(u5_mult_82_SUMB_36__10_) );
  FA_X1 u5_mult_82_S2_36_9 ( .A(u5_mult_82_ab_36__9_), .B(
        u5_mult_82_CARRYB_35__9_), .CI(u5_mult_82_SUMB_35__10_), .CO(
        u5_mult_82_CARRYB_36__9_), .S(u5_mult_82_SUMB_36__9_) );
  FA_X1 u5_mult_82_S2_36_8 ( .A(u5_mult_82_ab_36__8_), .B(
        u5_mult_82_CARRYB_35__8_), .CI(u5_mult_82_SUMB_35__9_), .CO(
        u5_mult_82_CARRYB_36__8_), .S(u5_mult_82_SUMB_36__8_) );
  FA_X1 u5_mult_82_S2_36_7 ( .A(u5_mult_82_ab_36__7_), .B(
        u5_mult_82_CARRYB_35__7_), .CI(u5_mult_82_SUMB_35__8_), .CO(
        u5_mult_82_CARRYB_36__7_), .S(u5_mult_82_SUMB_36__7_) );
  FA_X1 u5_mult_82_S2_36_6 ( .A(u5_mult_82_ab_36__6_), .B(
        u5_mult_82_CARRYB_35__6_), .CI(u5_mult_82_SUMB_35__7_), .CO(
        u5_mult_82_CARRYB_36__6_), .S(u5_mult_82_SUMB_36__6_) );
  FA_X1 u5_mult_82_S2_36_5 ( .A(u5_mult_82_ab_36__5_), .B(
        u5_mult_82_CARRYB_35__5_), .CI(u5_mult_82_SUMB_35__6_), .CO(
        u5_mult_82_CARRYB_36__5_), .S(u5_mult_82_SUMB_36__5_) );
  FA_X1 u5_mult_82_S2_36_4 ( .A(u5_mult_82_ab_36__4_), .B(
        u5_mult_82_CARRYB_35__4_), .CI(u5_mult_82_SUMB_35__5_), .CO(
        u5_mult_82_CARRYB_36__4_), .S(u5_mult_82_SUMB_36__4_) );
  FA_X1 u5_mult_82_S2_36_3 ( .A(u5_mult_82_ab_36__3_), .B(
        u5_mult_82_CARRYB_35__3_), .CI(u5_mult_82_SUMB_35__4_), .CO(
        u5_mult_82_CARRYB_36__3_), .S(u5_mult_82_SUMB_36__3_) );
  FA_X1 u5_mult_82_S2_36_2 ( .A(u5_mult_82_ab_36__2_), .B(
        u5_mult_82_CARRYB_35__2_), .CI(u5_mult_82_SUMB_35__3_), .CO(
        u5_mult_82_CARRYB_36__2_), .S(u5_mult_82_SUMB_36__2_) );
  FA_X1 u5_mult_82_S2_36_1 ( .A(u5_mult_82_ab_36__1_), .B(
        u5_mult_82_CARRYB_35__1_), .CI(u5_mult_82_SUMB_35__2_), .CO(
        u5_mult_82_CARRYB_36__1_), .S(u5_mult_82_SUMB_36__1_) );
  FA_X1 u5_mult_82_S1_36_0 ( .A(u5_mult_82_ab_36__0_), .B(
        u5_mult_82_CARRYB_35__0_), .CI(u5_mult_82_SUMB_35__1_), .CO(
        u5_mult_82_CARRYB_36__0_), .S(u5_N36) );
  FA_X1 u5_mult_82_S3_37_51 ( .A(u5_mult_82_ab_37__51_), .B(
        u5_mult_82_CARRYB_36__51_), .CI(u5_mult_82_ab_36__52_), .CO(
        u5_mult_82_CARRYB_37__51_), .S(u5_mult_82_SUMB_37__51_) );
  FA_X1 u5_mult_82_S2_37_50 ( .A(u5_mult_82_ab_37__50_), .B(
        u5_mult_82_CARRYB_36__50_), .CI(u5_mult_82_SUMB_36__51_), .CO(
        u5_mult_82_CARRYB_37__50_), .S(u5_mult_82_SUMB_37__50_) );
  FA_X1 u5_mult_82_S2_37_49 ( .A(u5_mult_82_ab_37__49_), .B(
        u5_mult_82_CARRYB_36__49_), .CI(u5_mult_82_SUMB_36__50_), .CO(
        u5_mult_82_CARRYB_37__49_), .S(u5_mult_82_SUMB_37__49_) );
  FA_X1 u5_mult_82_S2_37_48 ( .A(u5_mult_82_ab_37__48_), .B(
        u5_mult_82_CARRYB_36__48_), .CI(u5_mult_82_SUMB_36__49_), .CO(
        u5_mult_82_CARRYB_37__48_), .S(u5_mult_82_SUMB_37__48_) );
  FA_X1 u5_mult_82_S2_37_47 ( .A(u5_mult_82_ab_37__47_), .B(
        u5_mult_82_CARRYB_36__47_), .CI(u5_mult_82_SUMB_36__48_), .CO(
        u5_mult_82_CARRYB_37__47_), .S(u5_mult_82_SUMB_37__47_) );
  FA_X1 u5_mult_82_S2_37_46 ( .A(u5_mult_82_ab_37__46_), .B(
        u5_mult_82_CARRYB_36__46_), .CI(u5_mult_82_SUMB_36__47_), .CO(
        u5_mult_82_CARRYB_37__46_), .S(u5_mult_82_SUMB_37__46_) );
  FA_X1 u5_mult_82_S2_37_45 ( .A(u5_mult_82_ab_37__45_), .B(
        u5_mult_82_CARRYB_36__45_), .CI(u5_mult_82_SUMB_36__46_), .CO(
        u5_mult_82_CARRYB_37__45_), .S(u5_mult_82_SUMB_37__45_) );
  FA_X1 u5_mult_82_S2_37_44 ( .A(u5_mult_82_ab_37__44_), .B(
        u5_mult_82_CARRYB_36__44_), .CI(u5_mult_82_SUMB_36__45_), .CO(
        u5_mult_82_CARRYB_37__44_), .S(u5_mult_82_SUMB_37__44_) );
  FA_X1 u5_mult_82_S2_37_43 ( .A(u5_mult_82_ab_37__43_), .B(
        u5_mult_82_CARRYB_36__43_), .CI(u5_mult_82_SUMB_36__44_), .CO(
        u5_mult_82_CARRYB_37__43_), .S(u5_mult_82_SUMB_37__43_) );
  FA_X1 u5_mult_82_S2_37_42 ( .A(u5_mult_82_ab_37__42_), .B(
        u5_mult_82_CARRYB_36__42_), .CI(u5_mult_82_SUMB_36__43_), .CO(
        u5_mult_82_CARRYB_37__42_), .S(u5_mult_82_SUMB_37__42_) );
  FA_X1 u5_mult_82_S2_37_41 ( .A(u5_mult_82_ab_37__41_), .B(
        u5_mult_82_CARRYB_36__41_), .CI(u5_mult_82_SUMB_36__42_), .CO(
        u5_mult_82_CARRYB_37__41_), .S(u5_mult_82_SUMB_37__41_) );
  FA_X1 u5_mult_82_S2_37_40 ( .A(u5_mult_82_ab_37__40_), .B(
        u5_mult_82_CARRYB_36__40_), .CI(u5_mult_82_SUMB_36__41_), .CO(
        u5_mult_82_CARRYB_37__40_), .S(u5_mult_82_SUMB_37__40_) );
  FA_X1 u5_mult_82_S2_37_39 ( .A(u5_mult_82_ab_37__39_), .B(
        u5_mult_82_CARRYB_36__39_), .CI(u5_mult_82_SUMB_36__40_), .CO(
        u5_mult_82_CARRYB_37__39_), .S(u5_mult_82_SUMB_37__39_) );
  FA_X1 u5_mult_82_S2_37_38 ( .A(u5_mult_82_ab_37__38_), .B(
        u5_mult_82_CARRYB_36__38_), .CI(u5_mult_82_SUMB_36__39_), .CO(
        u5_mult_82_CARRYB_37__38_), .S(u5_mult_82_SUMB_37__38_) );
  FA_X1 u5_mult_82_S2_37_37 ( .A(u5_mult_82_ab_37__37_), .B(
        u5_mult_82_CARRYB_36__37_), .CI(u5_mult_82_SUMB_36__38_), .CO(
        u5_mult_82_CARRYB_37__37_), .S(u5_mult_82_SUMB_37__37_) );
  FA_X1 u5_mult_82_S2_37_36 ( .A(u5_mult_82_ab_37__36_), .B(
        u5_mult_82_CARRYB_36__36_), .CI(u5_mult_82_SUMB_36__37_), .CO(
        u5_mult_82_CARRYB_37__36_), .S(u5_mult_82_SUMB_37__36_) );
  FA_X1 u5_mult_82_S2_37_35 ( .A(u5_mult_82_ab_37__35_), .B(
        u5_mult_82_CARRYB_36__35_), .CI(u5_mult_82_SUMB_36__36_), .CO(
        u5_mult_82_CARRYB_37__35_), .S(u5_mult_82_SUMB_37__35_) );
  FA_X1 u5_mult_82_S2_37_34 ( .A(u5_mult_82_ab_37__34_), .B(
        u5_mult_82_CARRYB_36__34_), .CI(u5_mult_82_SUMB_36__35_), .CO(
        u5_mult_82_CARRYB_37__34_), .S(u5_mult_82_SUMB_37__34_) );
  FA_X1 u5_mult_82_S2_37_33 ( .A(u5_mult_82_ab_37__33_), .B(
        u5_mult_82_CARRYB_36__33_), .CI(u5_mult_82_SUMB_36__34_), .CO(
        u5_mult_82_CARRYB_37__33_), .S(u5_mult_82_SUMB_37__33_) );
  FA_X1 u5_mult_82_S2_37_32 ( .A(u5_mult_82_ab_37__32_), .B(
        u5_mult_82_CARRYB_36__32_), .CI(u5_mult_82_SUMB_36__33_), .CO(
        u5_mult_82_CARRYB_37__32_), .S(u5_mult_82_SUMB_37__32_) );
  FA_X1 u5_mult_82_S2_37_31 ( .A(u5_mult_82_ab_37__31_), .B(
        u5_mult_82_CARRYB_36__31_), .CI(u5_mult_82_SUMB_36__32_), .CO(
        u5_mult_82_CARRYB_37__31_), .S(u5_mult_82_SUMB_37__31_) );
  FA_X1 u5_mult_82_S2_37_30 ( .A(u5_mult_82_ab_37__30_), .B(
        u5_mult_82_CARRYB_36__30_), .CI(u5_mult_82_SUMB_36__31_), .CO(
        u5_mult_82_CARRYB_37__30_), .S(u5_mult_82_SUMB_37__30_) );
  FA_X1 u5_mult_82_S2_37_29 ( .A(u5_mult_82_ab_37__29_), .B(
        u5_mult_82_CARRYB_36__29_), .CI(u5_mult_82_SUMB_36__30_), .CO(
        u5_mult_82_CARRYB_37__29_), .S(u5_mult_82_SUMB_37__29_) );
  FA_X1 u5_mult_82_S2_37_28 ( .A(u5_mult_82_ab_37__28_), .B(
        u5_mult_82_CARRYB_36__28_), .CI(u5_mult_82_SUMB_36__29_), .CO(
        u5_mult_82_CARRYB_37__28_), .S(u5_mult_82_SUMB_37__28_) );
  FA_X1 u5_mult_82_S2_37_27 ( .A(u5_mult_82_ab_37__27_), .B(
        u5_mult_82_CARRYB_36__27_), .CI(u5_mult_82_SUMB_36__28_), .CO(
        u5_mult_82_CARRYB_37__27_), .S(u5_mult_82_SUMB_37__27_) );
  FA_X1 u5_mult_82_S2_37_26 ( .A(u5_mult_82_ab_37__26_), .B(
        u5_mult_82_CARRYB_36__26_), .CI(u5_mult_82_SUMB_36__27_), .CO(
        u5_mult_82_CARRYB_37__26_), .S(u5_mult_82_SUMB_37__26_) );
  FA_X1 u5_mult_82_S2_37_25 ( .A(u5_mult_82_ab_37__25_), .B(
        u5_mult_82_CARRYB_36__25_), .CI(u5_mult_82_SUMB_36__26_), .CO(
        u5_mult_82_CARRYB_37__25_), .S(u5_mult_82_SUMB_37__25_) );
  FA_X1 u5_mult_82_S2_37_24 ( .A(u5_mult_82_ab_37__24_), .B(
        u5_mult_82_CARRYB_36__24_), .CI(u5_mult_82_SUMB_36__25_), .CO(
        u5_mult_82_CARRYB_37__24_), .S(u5_mult_82_SUMB_37__24_) );
  FA_X1 u5_mult_82_S2_37_23 ( .A(u5_mult_82_ab_37__23_), .B(
        u5_mult_82_CARRYB_36__23_), .CI(u5_mult_82_SUMB_36__24_), .CO(
        u5_mult_82_CARRYB_37__23_), .S(u5_mult_82_SUMB_37__23_) );
  FA_X1 u5_mult_82_S2_37_22 ( .A(u5_mult_82_ab_37__22_), .B(
        u5_mult_82_CARRYB_36__22_), .CI(u5_mult_82_SUMB_36__23_), .CO(
        u5_mult_82_CARRYB_37__22_), .S(u5_mult_82_SUMB_37__22_) );
  FA_X1 u5_mult_82_S2_37_21 ( .A(u5_mult_82_ab_37__21_), .B(
        u5_mult_82_CARRYB_36__21_), .CI(u5_mult_82_SUMB_36__22_), .CO(
        u5_mult_82_CARRYB_37__21_), .S(u5_mult_82_SUMB_37__21_) );
  FA_X1 u5_mult_82_S2_37_20 ( .A(u5_mult_82_ab_37__20_), .B(
        u5_mult_82_CARRYB_36__20_), .CI(u5_mult_82_SUMB_36__21_), .CO(
        u5_mult_82_CARRYB_37__20_), .S(u5_mult_82_SUMB_37__20_) );
  FA_X1 u5_mult_82_S2_37_19 ( .A(u5_mult_82_ab_37__19_), .B(
        u5_mult_82_CARRYB_36__19_), .CI(u5_mult_82_SUMB_36__20_), .CO(
        u5_mult_82_CARRYB_37__19_), .S(u5_mult_82_SUMB_37__19_) );
  FA_X1 u5_mult_82_S2_37_18 ( .A(u5_mult_82_ab_37__18_), .B(
        u5_mult_82_CARRYB_36__18_), .CI(u5_mult_82_SUMB_36__19_), .CO(
        u5_mult_82_CARRYB_37__18_), .S(u5_mult_82_SUMB_37__18_) );
  FA_X1 u5_mult_82_S2_37_17 ( .A(u5_mult_82_ab_37__17_), .B(
        u5_mult_82_CARRYB_36__17_), .CI(u5_mult_82_SUMB_36__18_), .CO(
        u5_mult_82_CARRYB_37__17_), .S(u5_mult_82_SUMB_37__17_) );
  FA_X1 u5_mult_82_S2_37_16 ( .A(u5_mult_82_ab_37__16_), .B(
        u5_mult_82_CARRYB_36__16_), .CI(u5_mult_82_SUMB_36__17_), .CO(
        u5_mult_82_CARRYB_37__16_), .S(u5_mult_82_SUMB_37__16_) );
  FA_X1 u5_mult_82_S2_37_15 ( .A(u5_mult_82_ab_37__15_), .B(
        u5_mult_82_CARRYB_36__15_), .CI(u5_mult_82_SUMB_36__16_), .CO(
        u5_mult_82_CARRYB_37__15_), .S(u5_mult_82_SUMB_37__15_) );
  FA_X1 u5_mult_82_S2_37_14 ( .A(u5_mult_82_ab_37__14_), .B(
        u5_mult_82_CARRYB_36__14_), .CI(u5_mult_82_SUMB_36__15_), .CO(
        u5_mult_82_CARRYB_37__14_), .S(u5_mult_82_SUMB_37__14_) );
  FA_X1 u5_mult_82_S2_37_13 ( .A(u5_mult_82_ab_37__13_), .B(
        u5_mult_82_CARRYB_36__13_), .CI(u5_mult_82_SUMB_36__14_), .CO(
        u5_mult_82_CARRYB_37__13_), .S(u5_mult_82_SUMB_37__13_) );
  FA_X1 u5_mult_82_S2_37_12 ( .A(u5_mult_82_ab_37__12_), .B(
        u5_mult_82_CARRYB_36__12_), .CI(u5_mult_82_SUMB_36__13_), .CO(
        u5_mult_82_CARRYB_37__12_), .S(u5_mult_82_SUMB_37__12_) );
  FA_X1 u5_mult_82_S2_37_11 ( .A(u5_mult_82_ab_37__11_), .B(
        u5_mult_82_CARRYB_36__11_), .CI(u5_mult_82_SUMB_36__12_), .CO(
        u5_mult_82_CARRYB_37__11_), .S(u5_mult_82_SUMB_37__11_) );
  FA_X1 u5_mult_82_S2_37_10 ( .A(u5_mult_82_ab_37__10_), .B(
        u5_mult_82_CARRYB_36__10_), .CI(u5_mult_82_SUMB_36__11_), .CO(
        u5_mult_82_CARRYB_37__10_), .S(u5_mult_82_SUMB_37__10_) );
  FA_X1 u5_mult_82_S2_37_9 ( .A(u5_mult_82_ab_37__9_), .B(
        u5_mult_82_CARRYB_36__9_), .CI(u5_mult_82_SUMB_36__10_), .CO(
        u5_mult_82_CARRYB_37__9_), .S(u5_mult_82_SUMB_37__9_) );
  FA_X1 u5_mult_82_S2_37_8 ( .A(u5_mult_82_ab_37__8_), .B(
        u5_mult_82_CARRYB_36__8_), .CI(u5_mult_82_SUMB_36__9_), .CO(
        u5_mult_82_CARRYB_37__8_), .S(u5_mult_82_SUMB_37__8_) );
  FA_X1 u5_mult_82_S2_37_7 ( .A(u5_mult_82_ab_37__7_), .B(
        u5_mult_82_CARRYB_36__7_), .CI(u5_mult_82_SUMB_36__8_), .CO(
        u5_mult_82_CARRYB_37__7_), .S(u5_mult_82_SUMB_37__7_) );
  FA_X1 u5_mult_82_S2_37_6 ( .A(u5_mult_82_ab_37__6_), .B(
        u5_mult_82_CARRYB_36__6_), .CI(u5_mult_82_SUMB_36__7_), .CO(
        u5_mult_82_CARRYB_37__6_), .S(u5_mult_82_SUMB_37__6_) );
  FA_X1 u5_mult_82_S2_37_5 ( .A(u5_mult_82_ab_37__5_), .B(
        u5_mult_82_CARRYB_36__5_), .CI(u5_mult_82_SUMB_36__6_), .CO(
        u5_mult_82_CARRYB_37__5_), .S(u5_mult_82_SUMB_37__5_) );
  FA_X1 u5_mult_82_S2_37_4 ( .A(u5_mult_82_ab_37__4_), .B(
        u5_mult_82_CARRYB_36__4_), .CI(u5_mult_82_SUMB_36__5_), .CO(
        u5_mult_82_CARRYB_37__4_), .S(u5_mult_82_SUMB_37__4_) );
  FA_X1 u5_mult_82_S2_37_3 ( .A(u5_mult_82_ab_37__3_), .B(
        u5_mult_82_CARRYB_36__3_), .CI(u5_mult_82_SUMB_36__4_), .CO(
        u5_mult_82_CARRYB_37__3_), .S(u5_mult_82_SUMB_37__3_) );
  FA_X1 u5_mult_82_S2_37_2 ( .A(u5_mult_82_ab_37__2_), .B(
        u5_mult_82_CARRYB_36__2_), .CI(u5_mult_82_SUMB_36__3_), .CO(
        u5_mult_82_CARRYB_37__2_), .S(u5_mult_82_SUMB_37__2_) );
  FA_X1 u5_mult_82_S2_37_1 ( .A(u5_mult_82_ab_37__1_), .B(
        u5_mult_82_CARRYB_36__1_), .CI(u5_mult_82_SUMB_36__2_), .CO(
        u5_mult_82_CARRYB_37__1_), .S(u5_mult_82_SUMB_37__1_) );
  FA_X1 u5_mult_82_S1_37_0 ( .A(u5_mult_82_ab_37__0_), .B(
        u5_mult_82_CARRYB_36__0_), .CI(u5_mult_82_SUMB_36__1_), .CO(
        u5_mult_82_CARRYB_37__0_), .S(u5_N37) );
  FA_X1 u5_mult_82_S3_38_51 ( .A(u5_mult_82_ab_38__51_), .B(
        u5_mult_82_CARRYB_37__51_), .CI(u5_mult_82_ab_37__52_), .CO(
        u5_mult_82_CARRYB_38__51_), .S(u5_mult_82_SUMB_38__51_) );
  FA_X1 u5_mult_82_S2_38_50 ( .A(u5_mult_82_ab_38__50_), .B(
        u5_mult_82_CARRYB_37__50_), .CI(u5_mult_82_SUMB_37__51_), .CO(
        u5_mult_82_CARRYB_38__50_), .S(u5_mult_82_SUMB_38__50_) );
  FA_X1 u5_mult_82_S2_38_49 ( .A(u5_mult_82_ab_38__49_), .B(
        u5_mult_82_CARRYB_37__49_), .CI(u5_mult_82_SUMB_37__50_), .CO(
        u5_mult_82_CARRYB_38__49_), .S(u5_mult_82_SUMB_38__49_) );
  FA_X1 u5_mult_82_S2_38_48 ( .A(u5_mult_82_ab_38__48_), .B(
        u5_mult_82_CARRYB_37__48_), .CI(u5_mult_82_SUMB_37__49_), .CO(
        u5_mult_82_CARRYB_38__48_), .S(u5_mult_82_SUMB_38__48_) );
  FA_X1 u5_mult_82_S2_38_47 ( .A(u5_mult_82_ab_38__47_), .B(
        u5_mult_82_CARRYB_37__47_), .CI(u5_mult_82_SUMB_37__48_), .CO(
        u5_mult_82_CARRYB_38__47_), .S(u5_mult_82_SUMB_38__47_) );
  FA_X1 u5_mult_82_S2_38_46 ( .A(u5_mult_82_ab_38__46_), .B(
        u5_mult_82_CARRYB_37__46_), .CI(u5_mult_82_SUMB_37__47_), .CO(
        u5_mult_82_CARRYB_38__46_), .S(u5_mult_82_SUMB_38__46_) );
  FA_X1 u5_mult_82_S2_38_45 ( .A(u5_mult_82_ab_38__45_), .B(
        u5_mult_82_CARRYB_37__45_), .CI(u5_mult_82_SUMB_37__46_), .CO(
        u5_mult_82_CARRYB_38__45_), .S(u5_mult_82_SUMB_38__45_) );
  FA_X1 u5_mult_82_S2_38_44 ( .A(u5_mult_82_ab_38__44_), .B(
        u5_mult_82_CARRYB_37__44_), .CI(u5_mult_82_SUMB_37__45_), .CO(
        u5_mult_82_CARRYB_38__44_), .S(u5_mult_82_SUMB_38__44_) );
  FA_X1 u5_mult_82_S2_38_43 ( .A(u5_mult_82_ab_38__43_), .B(
        u5_mult_82_CARRYB_37__43_), .CI(u5_mult_82_SUMB_37__44_), .CO(
        u5_mult_82_CARRYB_38__43_), .S(u5_mult_82_SUMB_38__43_) );
  FA_X1 u5_mult_82_S2_38_42 ( .A(u5_mult_82_ab_38__42_), .B(
        u5_mult_82_CARRYB_37__42_), .CI(u5_mult_82_SUMB_37__43_), .CO(
        u5_mult_82_CARRYB_38__42_), .S(u5_mult_82_SUMB_38__42_) );
  FA_X1 u5_mult_82_S2_38_41 ( .A(u5_mult_82_ab_38__41_), .B(
        u5_mult_82_CARRYB_37__41_), .CI(u5_mult_82_SUMB_37__42_), .CO(
        u5_mult_82_CARRYB_38__41_), .S(u5_mult_82_SUMB_38__41_) );
  FA_X1 u5_mult_82_S2_38_40 ( .A(u5_mult_82_ab_38__40_), .B(
        u5_mult_82_CARRYB_37__40_), .CI(u5_mult_82_SUMB_37__41_), .CO(
        u5_mult_82_CARRYB_38__40_), .S(u5_mult_82_SUMB_38__40_) );
  FA_X1 u5_mult_82_S2_38_39 ( .A(u5_mult_82_ab_38__39_), .B(
        u5_mult_82_CARRYB_37__39_), .CI(u5_mult_82_SUMB_37__40_), .CO(
        u5_mult_82_CARRYB_38__39_), .S(u5_mult_82_SUMB_38__39_) );
  FA_X1 u5_mult_82_S2_38_38 ( .A(u5_mult_82_ab_38__38_), .B(
        u5_mult_82_CARRYB_37__38_), .CI(u5_mult_82_SUMB_37__39_), .CO(
        u5_mult_82_CARRYB_38__38_), .S(u5_mult_82_SUMB_38__38_) );
  FA_X1 u5_mult_82_S2_38_37 ( .A(u5_mult_82_ab_38__37_), .B(
        u5_mult_82_CARRYB_37__37_), .CI(u5_mult_82_SUMB_37__38_), .CO(
        u5_mult_82_CARRYB_38__37_), .S(u5_mult_82_SUMB_38__37_) );
  FA_X1 u5_mult_82_S2_38_36 ( .A(u5_mult_82_ab_38__36_), .B(
        u5_mult_82_CARRYB_37__36_), .CI(u5_mult_82_SUMB_37__37_), .CO(
        u5_mult_82_CARRYB_38__36_), .S(u5_mult_82_SUMB_38__36_) );
  FA_X1 u5_mult_82_S2_38_35 ( .A(u5_mult_82_ab_38__35_), .B(
        u5_mult_82_CARRYB_37__35_), .CI(u5_mult_82_SUMB_37__36_), .CO(
        u5_mult_82_CARRYB_38__35_), .S(u5_mult_82_SUMB_38__35_) );
  FA_X1 u5_mult_82_S2_38_34 ( .A(u5_mult_82_ab_38__34_), .B(
        u5_mult_82_CARRYB_37__34_), .CI(u5_mult_82_SUMB_37__35_), .CO(
        u5_mult_82_CARRYB_38__34_), .S(u5_mult_82_SUMB_38__34_) );
  FA_X1 u5_mult_82_S2_38_33 ( .A(u5_mult_82_ab_38__33_), .B(
        u5_mult_82_CARRYB_37__33_), .CI(u5_mult_82_SUMB_37__34_), .CO(
        u5_mult_82_CARRYB_38__33_), .S(u5_mult_82_SUMB_38__33_) );
  FA_X1 u5_mult_82_S2_38_32 ( .A(u5_mult_82_ab_38__32_), .B(
        u5_mult_82_CARRYB_37__32_), .CI(u5_mult_82_SUMB_37__33_), .CO(
        u5_mult_82_CARRYB_38__32_), .S(u5_mult_82_SUMB_38__32_) );
  FA_X1 u5_mult_82_S2_38_31 ( .A(u5_mult_82_ab_38__31_), .B(
        u5_mult_82_CARRYB_37__31_), .CI(u5_mult_82_SUMB_37__32_), .CO(
        u5_mult_82_CARRYB_38__31_), .S(u5_mult_82_SUMB_38__31_) );
  FA_X1 u5_mult_82_S2_38_30 ( .A(u5_mult_82_ab_38__30_), .B(
        u5_mult_82_CARRYB_37__30_), .CI(u5_mult_82_SUMB_37__31_), .CO(
        u5_mult_82_CARRYB_38__30_), .S(u5_mult_82_SUMB_38__30_) );
  FA_X1 u5_mult_82_S2_38_29 ( .A(u5_mult_82_ab_38__29_), .B(
        u5_mult_82_CARRYB_37__29_), .CI(u5_mult_82_SUMB_37__30_), .CO(
        u5_mult_82_CARRYB_38__29_), .S(u5_mult_82_SUMB_38__29_) );
  FA_X1 u5_mult_82_S2_38_28 ( .A(u5_mult_82_ab_38__28_), .B(
        u5_mult_82_CARRYB_37__28_), .CI(u5_mult_82_SUMB_37__29_), .CO(
        u5_mult_82_CARRYB_38__28_), .S(u5_mult_82_SUMB_38__28_) );
  FA_X1 u5_mult_82_S2_38_27 ( .A(u5_mult_82_ab_38__27_), .B(
        u5_mult_82_CARRYB_37__27_), .CI(u5_mult_82_SUMB_37__28_), .CO(
        u5_mult_82_CARRYB_38__27_), .S(u5_mult_82_SUMB_38__27_) );
  FA_X1 u5_mult_82_S2_38_26 ( .A(u5_mult_82_ab_38__26_), .B(
        u5_mult_82_CARRYB_37__26_), .CI(u5_mult_82_SUMB_37__27_), .CO(
        u5_mult_82_CARRYB_38__26_), .S(u5_mult_82_SUMB_38__26_) );
  FA_X1 u5_mult_82_S2_38_25 ( .A(u5_mult_82_ab_38__25_), .B(
        u5_mult_82_CARRYB_37__25_), .CI(u5_mult_82_SUMB_37__26_), .CO(
        u5_mult_82_CARRYB_38__25_), .S(u5_mult_82_SUMB_38__25_) );
  FA_X1 u5_mult_82_S2_38_24 ( .A(u5_mult_82_ab_38__24_), .B(
        u5_mult_82_CARRYB_37__24_), .CI(u5_mult_82_SUMB_37__25_), .CO(
        u5_mult_82_CARRYB_38__24_), .S(u5_mult_82_SUMB_38__24_) );
  FA_X1 u5_mult_82_S2_38_23 ( .A(u5_mult_82_ab_38__23_), .B(
        u5_mult_82_CARRYB_37__23_), .CI(u5_mult_82_SUMB_37__24_), .CO(
        u5_mult_82_CARRYB_38__23_), .S(u5_mult_82_SUMB_38__23_) );
  FA_X1 u5_mult_82_S2_38_22 ( .A(u5_mult_82_ab_38__22_), .B(
        u5_mult_82_CARRYB_37__22_), .CI(u5_mult_82_SUMB_37__23_), .CO(
        u5_mult_82_CARRYB_38__22_), .S(u5_mult_82_SUMB_38__22_) );
  FA_X1 u5_mult_82_S2_38_21 ( .A(u5_mult_82_ab_38__21_), .B(
        u5_mult_82_CARRYB_37__21_), .CI(u5_mult_82_SUMB_37__22_), .CO(
        u5_mult_82_CARRYB_38__21_), .S(u5_mult_82_SUMB_38__21_) );
  FA_X1 u5_mult_82_S2_38_20 ( .A(u5_mult_82_ab_38__20_), .B(
        u5_mult_82_CARRYB_37__20_), .CI(u5_mult_82_SUMB_37__21_), .CO(
        u5_mult_82_CARRYB_38__20_), .S(u5_mult_82_SUMB_38__20_) );
  FA_X1 u5_mult_82_S2_38_19 ( .A(u5_mult_82_ab_38__19_), .B(
        u5_mult_82_CARRYB_37__19_), .CI(u5_mult_82_SUMB_37__20_), .CO(
        u5_mult_82_CARRYB_38__19_), .S(u5_mult_82_SUMB_38__19_) );
  FA_X1 u5_mult_82_S2_38_18 ( .A(u5_mult_82_ab_38__18_), .B(
        u5_mult_82_CARRYB_37__18_), .CI(u5_mult_82_SUMB_37__19_), .CO(
        u5_mult_82_CARRYB_38__18_), .S(u5_mult_82_SUMB_38__18_) );
  FA_X1 u5_mult_82_S2_38_17 ( .A(u5_mult_82_ab_38__17_), .B(
        u5_mult_82_CARRYB_37__17_), .CI(u5_mult_82_SUMB_37__18_), .CO(
        u5_mult_82_CARRYB_38__17_), .S(u5_mult_82_SUMB_38__17_) );
  FA_X1 u5_mult_82_S2_38_16 ( .A(u5_mult_82_ab_38__16_), .B(
        u5_mult_82_CARRYB_37__16_), .CI(u5_mult_82_SUMB_37__17_), .CO(
        u5_mult_82_CARRYB_38__16_), .S(u5_mult_82_SUMB_38__16_) );
  FA_X1 u5_mult_82_S2_38_15 ( .A(u5_mult_82_ab_38__15_), .B(
        u5_mult_82_CARRYB_37__15_), .CI(u5_mult_82_SUMB_37__16_), .CO(
        u5_mult_82_CARRYB_38__15_), .S(u5_mult_82_SUMB_38__15_) );
  FA_X1 u5_mult_82_S2_38_14 ( .A(u5_mult_82_ab_38__14_), .B(
        u5_mult_82_CARRYB_37__14_), .CI(u5_mult_82_SUMB_37__15_), .CO(
        u5_mult_82_CARRYB_38__14_), .S(u5_mult_82_SUMB_38__14_) );
  FA_X1 u5_mult_82_S2_38_13 ( .A(u5_mult_82_ab_38__13_), .B(
        u5_mult_82_CARRYB_37__13_), .CI(u5_mult_82_SUMB_37__14_), .CO(
        u5_mult_82_CARRYB_38__13_), .S(u5_mult_82_SUMB_38__13_) );
  FA_X1 u5_mult_82_S2_38_12 ( .A(u5_mult_82_ab_38__12_), .B(
        u5_mult_82_CARRYB_37__12_), .CI(u5_mult_82_SUMB_37__13_), .CO(
        u5_mult_82_CARRYB_38__12_), .S(u5_mult_82_SUMB_38__12_) );
  FA_X1 u5_mult_82_S2_38_11 ( .A(u5_mult_82_ab_38__11_), .B(
        u5_mult_82_CARRYB_37__11_), .CI(u5_mult_82_SUMB_37__12_), .CO(
        u5_mult_82_CARRYB_38__11_), .S(u5_mult_82_SUMB_38__11_) );
  FA_X1 u5_mult_82_S2_38_10 ( .A(u5_mult_82_ab_38__10_), .B(
        u5_mult_82_CARRYB_37__10_), .CI(u5_mult_82_SUMB_37__11_), .CO(
        u5_mult_82_CARRYB_38__10_), .S(u5_mult_82_SUMB_38__10_) );
  FA_X1 u5_mult_82_S2_38_9 ( .A(u5_mult_82_ab_38__9_), .B(
        u5_mult_82_CARRYB_37__9_), .CI(u5_mult_82_SUMB_37__10_), .CO(
        u5_mult_82_CARRYB_38__9_), .S(u5_mult_82_SUMB_38__9_) );
  FA_X1 u5_mult_82_S2_38_8 ( .A(u5_mult_82_ab_38__8_), .B(
        u5_mult_82_CARRYB_37__8_), .CI(u5_mult_82_SUMB_37__9_), .CO(
        u5_mult_82_CARRYB_38__8_), .S(u5_mult_82_SUMB_38__8_) );
  FA_X1 u5_mult_82_S2_38_7 ( .A(u5_mult_82_ab_38__7_), .B(
        u5_mult_82_CARRYB_37__7_), .CI(u5_mult_82_SUMB_37__8_), .CO(
        u5_mult_82_CARRYB_38__7_), .S(u5_mult_82_SUMB_38__7_) );
  FA_X1 u5_mult_82_S2_38_6 ( .A(u5_mult_82_ab_38__6_), .B(
        u5_mult_82_CARRYB_37__6_), .CI(u5_mult_82_SUMB_37__7_), .CO(
        u5_mult_82_CARRYB_38__6_), .S(u5_mult_82_SUMB_38__6_) );
  FA_X1 u5_mult_82_S2_38_5 ( .A(u5_mult_82_ab_38__5_), .B(
        u5_mult_82_CARRYB_37__5_), .CI(u5_mult_82_SUMB_37__6_), .CO(
        u5_mult_82_CARRYB_38__5_), .S(u5_mult_82_SUMB_38__5_) );
  FA_X1 u5_mult_82_S2_38_4 ( .A(u5_mult_82_ab_38__4_), .B(
        u5_mult_82_CARRYB_37__4_), .CI(u5_mult_82_SUMB_37__5_), .CO(
        u5_mult_82_CARRYB_38__4_), .S(u5_mult_82_SUMB_38__4_) );
  FA_X1 u5_mult_82_S2_38_3 ( .A(u5_mult_82_ab_38__3_), .B(
        u5_mult_82_CARRYB_37__3_), .CI(u5_mult_82_SUMB_37__4_), .CO(
        u5_mult_82_CARRYB_38__3_), .S(u5_mult_82_SUMB_38__3_) );
  FA_X1 u5_mult_82_S2_38_2 ( .A(u5_mult_82_ab_38__2_), .B(
        u5_mult_82_CARRYB_37__2_), .CI(u5_mult_82_SUMB_37__3_), .CO(
        u5_mult_82_CARRYB_38__2_), .S(u5_mult_82_SUMB_38__2_) );
  FA_X1 u5_mult_82_S2_38_1 ( .A(u5_mult_82_ab_38__1_), .B(
        u5_mult_82_CARRYB_37__1_), .CI(u5_mult_82_SUMB_37__2_), .CO(
        u5_mult_82_CARRYB_38__1_), .S(u5_mult_82_SUMB_38__1_) );
  FA_X1 u5_mult_82_S1_38_0 ( .A(u5_mult_82_ab_38__0_), .B(
        u5_mult_82_CARRYB_37__0_), .CI(u5_mult_82_SUMB_37__1_), .CO(
        u5_mult_82_CARRYB_38__0_), .S(u5_N38) );
  FA_X1 u5_mult_82_S3_39_51 ( .A(u5_mult_82_ab_39__51_), .B(
        u5_mult_82_CARRYB_38__51_), .CI(u5_mult_82_ab_38__52_), .CO(
        u5_mult_82_CARRYB_39__51_), .S(u5_mult_82_SUMB_39__51_) );
  FA_X1 u5_mult_82_S2_39_50 ( .A(u5_mult_82_ab_39__50_), .B(
        u5_mult_82_CARRYB_38__50_), .CI(u5_mult_82_SUMB_38__51_), .CO(
        u5_mult_82_CARRYB_39__50_), .S(u5_mult_82_SUMB_39__50_) );
  FA_X1 u5_mult_82_S2_39_49 ( .A(u5_mult_82_ab_39__49_), .B(
        u5_mult_82_CARRYB_38__49_), .CI(u5_mult_82_SUMB_38__50_), .CO(
        u5_mult_82_CARRYB_39__49_), .S(u5_mult_82_SUMB_39__49_) );
  FA_X1 u5_mult_82_S2_39_48 ( .A(u5_mult_82_ab_39__48_), .B(
        u5_mult_82_CARRYB_38__48_), .CI(u5_mult_82_SUMB_38__49_), .CO(
        u5_mult_82_CARRYB_39__48_), .S(u5_mult_82_SUMB_39__48_) );
  FA_X1 u5_mult_82_S2_39_47 ( .A(u5_mult_82_ab_39__47_), .B(
        u5_mult_82_CARRYB_38__47_), .CI(u5_mult_82_SUMB_38__48_), .CO(
        u5_mult_82_CARRYB_39__47_), .S(u5_mult_82_SUMB_39__47_) );
  FA_X1 u5_mult_82_S2_39_46 ( .A(u5_mult_82_ab_39__46_), .B(
        u5_mult_82_CARRYB_38__46_), .CI(u5_mult_82_SUMB_38__47_), .CO(
        u5_mult_82_CARRYB_39__46_), .S(u5_mult_82_SUMB_39__46_) );
  FA_X1 u5_mult_82_S2_39_45 ( .A(u5_mult_82_ab_39__45_), .B(
        u5_mult_82_CARRYB_38__45_), .CI(u5_mult_82_SUMB_38__46_), .CO(
        u5_mult_82_CARRYB_39__45_), .S(u5_mult_82_SUMB_39__45_) );
  FA_X1 u5_mult_82_S2_39_44 ( .A(u5_mult_82_ab_39__44_), .B(
        u5_mult_82_CARRYB_38__44_), .CI(u5_mult_82_SUMB_38__45_), .CO(
        u5_mult_82_CARRYB_39__44_), .S(u5_mult_82_SUMB_39__44_) );
  FA_X1 u5_mult_82_S2_39_43 ( .A(u5_mult_82_ab_39__43_), .B(
        u5_mult_82_CARRYB_38__43_), .CI(u5_mult_82_SUMB_38__44_), .CO(
        u5_mult_82_CARRYB_39__43_), .S(u5_mult_82_SUMB_39__43_) );
  FA_X1 u5_mult_82_S2_39_42 ( .A(u5_mult_82_ab_39__42_), .B(
        u5_mult_82_CARRYB_38__42_), .CI(u5_mult_82_SUMB_38__43_), .CO(
        u5_mult_82_CARRYB_39__42_), .S(u5_mult_82_SUMB_39__42_) );
  FA_X1 u5_mult_82_S2_39_41 ( .A(u5_mult_82_ab_39__41_), .B(
        u5_mult_82_CARRYB_38__41_), .CI(u5_mult_82_SUMB_38__42_), .CO(
        u5_mult_82_CARRYB_39__41_), .S(u5_mult_82_SUMB_39__41_) );
  FA_X1 u5_mult_82_S2_39_40 ( .A(u5_mult_82_ab_39__40_), .B(
        u5_mult_82_CARRYB_38__40_), .CI(u5_mult_82_SUMB_38__41_), .CO(
        u5_mult_82_CARRYB_39__40_), .S(u5_mult_82_SUMB_39__40_) );
  FA_X1 u5_mult_82_S2_39_39 ( .A(u5_mult_82_ab_39__39_), .B(
        u5_mult_82_CARRYB_38__39_), .CI(u5_mult_82_SUMB_38__40_), .CO(
        u5_mult_82_CARRYB_39__39_), .S(u5_mult_82_SUMB_39__39_) );
  FA_X1 u5_mult_82_S2_39_38 ( .A(u5_mult_82_ab_39__38_), .B(
        u5_mult_82_CARRYB_38__38_), .CI(u5_mult_82_SUMB_38__39_), .CO(
        u5_mult_82_CARRYB_39__38_), .S(u5_mult_82_SUMB_39__38_) );
  FA_X1 u5_mult_82_S2_39_37 ( .A(u5_mult_82_ab_39__37_), .B(
        u5_mult_82_CARRYB_38__37_), .CI(u5_mult_82_SUMB_38__38_), .CO(
        u5_mult_82_CARRYB_39__37_), .S(u5_mult_82_SUMB_39__37_) );
  FA_X1 u5_mult_82_S2_39_36 ( .A(u5_mult_82_ab_39__36_), .B(
        u5_mult_82_CARRYB_38__36_), .CI(u5_mult_82_SUMB_38__37_), .CO(
        u5_mult_82_CARRYB_39__36_), .S(u5_mult_82_SUMB_39__36_) );
  FA_X1 u5_mult_82_S2_39_35 ( .A(u5_mult_82_ab_39__35_), .B(
        u5_mult_82_CARRYB_38__35_), .CI(u5_mult_82_SUMB_38__36_), .CO(
        u5_mult_82_CARRYB_39__35_), .S(u5_mult_82_SUMB_39__35_) );
  FA_X1 u5_mult_82_S2_39_34 ( .A(u5_mult_82_ab_39__34_), .B(
        u5_mult_82_CARRYB_38__34_), .CI(u5_mult_82_SUMB_38__35_), .CO(
        u5_mult_82_CARRYB_39__34_), .S(u5_mult_82_SUMB_39__34_) );
  FA_X1 u5_mult_82_S2_39_33 ( .A(u5_mult_82_ab_39__33_), .B(
        u5_mult_82_CARRYB_38__33_), .CI(u5_mult_82_SUMB_38__34_), .CO(
        u5_mult_82_CARRYB_39__33_), .S(u5_mult_82_SUMB_39__33_) );
  FA_X1 u5_mult_82_S2_39_32 ( .A(u5_mult_82_ab_39__32_), .B(
        u5_mult_82_CARRYB_38__32_), .CI(u5_mult_82_SUMB_38__33_), .CO(
        u5_mult_82_CARRYB_39__32_), .S(u5_mult_82_SUMB_39__32_) );
  FA_X1 u5_mult_82_S2_39_31 ( .A(u5_mult_82_ab_39__31_), .B(
        u5_mult_82_CARRYB_38__31_), .CI(u5_mult_82_SUMB_38__32_), .CO(
        u5_mult_82_CARRYB_39__31_), .S(u5_mult_82_SUMB_39__31_) );
  FA_X1 u5_mult_82_S2_39_30 ( .A(u5_mult_82_ab_39__30_), .B(
        u5_mult_82_CARRYB_38__30_), .CI(u5_mult_82_SUMB_38__31_), .CO(
        u5_mult_82_CARRYB_39__30_), .S(u5_mult_82_SUMB_39__30_) );
  FA_X1 u5_mult_82_S2_39_29 ( .A(u5_mult_82_ab_39__29_), .B(
        u5_mult_82_CARRYB_38__29_), .CI(u5_mult_82_SUMB_38__30_), .CO(
        u5_mult_82_CARRYB_39__29_), .S(u5_mult_82_SUMB_39__29_) );
  FA_X1 u5_mult_82_S2_39_28 ( .A(u5_mult_82_ab_39__28_), .B(
        u5_mult_82_CARRYB_38__28_), .CI(u5_mult_82_SUMB_38__29_), .CO(
        u5_mult_82_CARRYB_39__28_), .S(u5_mult_82_SUMB_39__28_) );
  FA_X1 u5_mult_82_S2_39_27 ( .A(u5_mult_82_ab_39__27_), .B(
        u5_mult_82_CARRYB_38__27_), .CI(u5_mult_82_SUMB_38__28_), .CO(
        u5_mult_82_CARRYB_39__27_), .S(u5_mult_82_SUMB_39__27_) );
  FA_X1 u5_mult_82_S2_39_26 ( .A(u5_mult_82_ab_39__26_), .B(
        u5_mult_82_CARRYB_38__26_), .CI(u5_mult_82_SUMB_38__27_), .CO(
        u5_mult_82_CARRYB_39__26_), .S(u5_mult_82_SUMB_39__26_) );
  FA_X1 u5_mult_82_S2_39_25 ( .A(u5_mult_82_ab_39__25_), .B(
        u5_mult_82_CARRYB_38__25_), .CI(u5_mult_82_SUMB_38__26_), .CO(
        u5_mult_82_CARRYB_39__25_), .S(u5_mult_82_SUMB_39__25_) );
  FA_X1 u5_mult_82_S2_39_24 ( .A(u5_mult_82_ab_39__24_), .B(
        u5_mult_82_CARRYB_38__24_), .CI(u5_mult_82_SUMB_38__25_), .CO(
        u5_mult_82_CARRYB_39__24_), .S(u5_mult_82_SUMB_39__24_) );
  FA_X1 u5_mult_82_S2_39_23 ( .A(u5_mult_82_ab_39__23_), .B(
        u5_mult_82_CARRYB_38__23_), .CI(u5_mult_82_SUMB_38__24_), .CO(
        u5_mult_82_CARRYB_39__23_), .S(u5_mult_82_SUMB_39__23_) );
  FA_X1 u5_mult_82_S2_39_22 ( .A(u5_mult_82_ab_39__22_), .B(
        u5_mult_82_CARRYB_38__22_), .CI(u5_mult_82_SUMB_38__23_), .CO(
        u5_mult_82_CARRYB_39__22_), .S(u5_mult_82_SUMB_39__22_) );
  FA_X1 u5_mult_82_S2_39_21 ( .A(u5_mult_82_ab_39__21_), .B(
        u5_mult_82_CARRYB_38__21_), .CI(u5_mult_82_SUMB_38__22_), .CO(
        u5_mult_82_CARRYB_39__21_), .S(u5_mult_82_SUMB_39__21_) );
  FA_X1 u5_mult_82_S2_39_20 ( .A(u5_mult_82_ab_39__20_), .B(
        u5_mult_82_CARRYB_38__20_), .CI(u5_mult_82_SUMB_38__21_), .CO(
        u5_mult_82_CARRYB_39__20_), .S(u5_mult_82_SUMB_39__20_) );
  FA_X1 u5_mult_82_S2_39_19 ( .A(u5_mult_82_ab_39__19_), .B(
        u5_mult_82_CARRYB_38__19_), .CI(u5_mult_82_SUMB_38__20_), .CO(
        u5_mult_82_CARRYB_39__19_), .S(u5_mult_82_SUMB_39__19_) );
  FA_X1 u5_mult_82_S2_39_18 ( .A(u5_mult_82_ab_39__18_), .B(
        u5_mult_82_CARRYB_38__18_), .CI(u5_mult_82_SUMB_38__19_), .CO(
        u5_mult_82_CARRYB_39__18_), .S(u5_mult_82_SUMB_39__18_) );
  FA_X1 u5_mult_82_S2_39_17 ( .A(u5_mult_82_ab_39__17_), .B(
        u5_mult_82_CARRYB_38__17_), .CI(u5_mult_82_SUMB_38__18_), .CO(
        u5_mult_82_CARRYB_39__17_), .S(u5_mult_82_SUMB_39__17_) );
  FA_X1 u5_mult_82_S2_39_16 ( .A(u5_mult_82_ab_39__16_), .B(
        u5_mult_82_CARRYB_38__16_), .CI(u5_mult_82_SUMB_38__17_), .CO(
        u5_mult_82_CARRYB_39__16_), .S(u5_mult_82_SUMB_39__16_) );
  FA_X1 u5_mult_82_S2_39_15 ( .A(u5_mult_82_ab_39__15_), .B(
        u5_mult_82_CARRYB_38__15_), .CI(u5_mult_82_SUMB_38__16_), .CO(
        u5_mult_82_CARRYB_39__15_), .S(u5_mult_82_SUMB_39__15_) );
  FA_X1 u5_mult_82_S2_39_14 ( .A(u5_mult_82_ab_39__14_), .B(
        u5_mult_82_CARRYB_38__14_), .CI(u5_mult_82_SUMB_38__15_), .CO(
        u5_mult_82_CARRYB_39__14_), .S(u5_mult_82_SUMB_39__14_) );
  FA_X1 u5_mult_82_S2_39_13 ( .A(u5_mult_82_ab_39__13_), .B(
        u5_mult_82_CARRYB_38__13_), .CI(u5_mult_82_SUMB_38__14_), .CO(
        u5_mult_82_CARRYB_39__13_), .S(u5_mult_82_SUMB_39__13_) );
  FA_X1 u5_mult_82_S2_39_12 ( .A(u5_mult_82_ab_39__12_), .B(
        u5_mult_82_CARRYB_38__12_), .CI(u5_mult_82_SUMB_38__13_), .CO(
        u5_mult_82_CARRYB_39__12_), .S(u5_mult_82_SUMB_39__12_) );
  FA_X1 u5_mult_82_S2_39_11 ( .A(u5_mult_82_ab_39__11_), .B(
        u5_mult_82_CARRYB_38__11_), .CI(u5_mult_82_SUMB_38__12_), .CO(
        u5_mult_82_CARRYB_39__11_), .S(u5_mult_82_SUMB_39__11_) );
  FA_X1 u5_mult_82_S2_39_10 ( .A(u5_mult_82_ab_39__10_), .B(
        u5_mult_82_CARRYB_38__10_), .CI(u5_mult_82_SUMB_38__11_), .CO(
        u5_mult_82_CARRYB_39__10_), .S(u5_mult_82_SUMB_39__10_) );
  FA_X1 u5_mult_82_S2_39_9 ( .A(u5_mult_82_ab_39__9_), .B(
        u5_mult_82_CARRYB_38__9_), .CI(u5_mult_82_SUMB_38__10_), .CO(
        u5_mult_82_CARRYB_39__9_), .S(u5_mult_82_SUMB_39__9_) );
  FA_X1 u5_mult_82_S2_39_8 ( .A(u5_mult_82_ab_39__8_), .B(
        u5_mult_82_CARRYB_38__8_), .CI(u5_mult_82_SUMB_38__9_), .CO(
        u5_mult_82_CARRYB_39__8_), .S(u5_mult_82_SUMB_39__8_) );
  FA_X1 u5_mult_82_S2_39_7 ( .A(u5_mult_82_ab_39__7_), .B(
        u5_mult_82_CARRYB_38__7_), .CI(u5_mult_82_SUMB_38__8_), .CO(
        u5_mult_82_CARRYB_39__7_), .S(u5_mult_82_SUMB_39__7_) );
  FA_X1 u5_mult_82_S2_39_6 ( .A(u5_mult_82_ab_39__6_), .B(
        u5_mult_82_CARRYB_38__6_), .CI(u5_mult_82_SUMB_38__7_), .CO(
        u5_mult_82_CARRYB_39__6_), .S(u5_mult_82_SUMB_39__6_) );
  FA_X1 u5_mult_82_S2_39_5 ( .A(u5_mult_82_ab_39__5_), .B(
        u5_mult_82_CARRYB_38__5_), .CI(u5_mult_82_SUMB_38__6_), .CO(
        u5_mult_82_CARRYB_39__5_), .S(u5_mult_82_SUMB_39__5_) );
  FA_X1 u5_mult_82_S2_39_4 ( .A(u5_mult_82_ab_39__4_), .B(
        u5_mult_82_CARRYB_38__4_), .CI(u5_mult_82_SUMB_38__5_), .CO(
        u5_mult_82_CARRYB_39__4_), .S(u5_mult_82_SUMB_39__4_) );
  FA_X1 u5_mult_82_S2_39_3 ( .A(u5_mult_82_ab_39__3_), .B(
        u5_mult_82_CARRYB_38__3_), .CI(u5_mult_82_SUMB_38__4_), .CO(
        u5_mult_82_CARRYB_39__3_), .S(u5_mult_82_SUMB_39__3_) );
  FA_X1 u5_mult_82_S2_39_2 ( .A(u5_mult_82_ab_39__2_), .B(
        u5_mult_82_CARRYB_38__2_), .CI(u5_mult_82_SUMB_38__3_), .CO(
        u5_mult_82_CARRYB_39__2_), .S(u5_mult_82_SUMB_39__2_) );
  FA_X1 u5_mult_82_S2_39_1 ( .A(u5_mult_82_ab_39__1_), .B(
        u5_mult_82_CARRYB_38__1_), .CI(u5_mult_82_SUMB_38__2_), .CO(
        u5_mult_82_CARRYB_39__1_), .S(u5_mult_82_SUMB_39__1_) );
  FA_X1 u5_mult_82_S1_39_0 ( .A(u5_mult_82_ab_39__0_), .B(
        u5_mult_82_CARRYB_38__0_), .CI(u5_mult_82_SUMB_38__1_), .CO(
        u5_mult_82_CARRYB_39__0_), .S(u5_N39) );
  FA_X1 u5_mult_82_S3_40_51 ( .A(u5_mult_82_ab_40__51_), .B(
        u5_mult_82_CARRYB_39__51_), .CI(u5_mult_82_ab_39__52_), .CO(
        u5_mult_82_CARRYB_40__51_), .S(u5_mult_82_SUMB_40__51_) );
  FA_X1 u5_mult_82_S2_40_50 ( .A(u5_mult_82_ab_40__50_), .B(
        u5_mult_82_CARRYB_39__50_), .CI(u5_mult_82_SUMB_39__51_), .CO(
        u5_mult_82_CARRYB_40__50_), .S(u5_mult_82_SUMB_40__50_) );
  FA_X1 u5_mult_82_S2_40_49 ( .A(u5_mult_82_ab_40__49_), .B(
        u5_mult_82_CARRYB_39__49_), .CI(u5_mult_82_SUMB_39__50_), .CO(
        u5_mult_82_CARRYB_40__49_), .S(u5_mult_82_SUMB_40__49_) );
  FA_X1 u5_mult_82_S2_40_48 ( .A(u5_mult_82_ab_40__48_), .B(
        u5_mult_82_CARRYB_39__48_), .CI(u5_mult_82_SUMB_39__49_), .CO(
        u5_mult_82_CARRYB_40__48_), .S(u5_mult_82_SUMB_40__48_) );
  FA_X1 u5_mult_82_S2_40_47 ( .A(u5_mult_82_ab_40__47_), .B(
        u5_mult_82_CARRYB_39__47_), .CI(u5_mult_82_SUMB_39__48_), .CO(
        u5_mult_82_CARRYB_40__47_), .S(u5_mult_82_SUMB_40__47_) );
  FA_X1 u5_mult_82_S2_40_46 ( .A(u5_mult_82_ab_40__46_), .B(
        u5_mult_82_CARRYB_39__46_), .CI(u5_mult_82_SUMB_39__47_), .CO(
        u5_mult_82_CARRYB_40__46_), .S(u5_mult_82_SUMB_40__46_) );
  FA_X1 u5_mult_82_S2_40_45 ( .A(u5_mult_82_ab_40__45_), .B(
        u5_mult_82_CARRYB_39__45_), .CI(u5_mult_82_SUMB_39__46_), .CO(
        u5_mult_82_CARRYB_40__45_), .S(u5_mult_82_SUMB_40__45_) );
  FA_X1 u5_mult_82_S2_40_44 ( .A(u5_mult_82_ab_40__44_), .B(
        u5_mult_82_CARRYB_39__44_), .CI(u5_mult_82_SUMB_39__45_), .CO(
        u5_mult_82_CARRYB_40__44_), .S(u5_mult_82_SUMB_40__44_) );
  FA_X1 u5_mult_82_S2_40_43 ( .A(u5_mult_82_ab_40__43_), .B(
        u5_mult_82_CARRYB_39__43_), .CI(u5_mult_82_SUMB_39__44_), .CO(
        u5_mult_82_CARRYB_40__43_), .S(u5_mult_82_SUMB_40__43_) );
  FA_X1 u5_mult_82_S2_40_42 ( .A(u5_mult_82_ab_40__42_), .B(
        u5_mult_82_CARRYB_39__42_), .CI(u5_mult_82_SUMB_39__43_), .CO(
        u5_mult_82_CARRYB_40__42_), .S(u5_mult_82_SUMB_40__42_) );
  FA_X1 u5_mult_82_S2_40_41 ( .A(u5_mult_82_ab_40__41_), .B(
        u5_mult_82_CARRYB_39__41_), .CI(u5_mult_82_SUMB_39__42_), .CO(
        u5_mult_82_CARRYB_40__41_), .S(u5_mult_82_SUMB_40__41_) );
  FA_X1 u5_mult_82_S2_40_40 ( .A(u5_mult_82_ab_40__40_), .B(
        u5_mult_82_CARRYB_39__40_), .CI(u5_mult_82_SUMB_39__41_), .CO(
        u5_mult_82_CARRYB_40__40_), .S(u5_mult_82_SUMB_40__40_) );
  FA_X1 u5_mult_82_S2_40_39 ( .A(u5_mult_82_ab_40__39_), .B(
        u5_mult_82_CARRYB_39__39_), .CI(u5_mult_82_SUMB_39__40_), .CO(
        u5_mult_82_CARRYB_40__39_), .S(u5_mult_82_SUMB_40__39_) );
  FA_X1 u5_mult_82_S2_40_38 ( .A(u5_mult_82_ab_40__38_), .B(
        u5_mult_82_CARRYB_39__38_), .CI(u5_mult_82_SUMB_39__39_), .CO(
        u5_mult_82_CARRYB_40__38_), .S(u5_mult_82_SUMB_40__38_) );
  FA_X1 u5_mult_82_S2_40_37 ( .A(u5_mult_82_ab_40__37_), .B(
        u5_mult_82_CARRYB_39__37_), .CI(u5_mult_82_SUMB_39__38_), .CO(
        u5_mult_82_CARRYB_40__37_), .S(u5_mult_82_SUMB_40__37_) );
  FA_X1 u5_mult_82_S2_40_36 ( .A(u5_mult_82_ab_40__36_), .B(
        u5_mult_82_CARRYB_39__36_), .CI(u5_mult_82_SUMB_39__37_), .CO(
        u5_mult_82_CARRYB_40__36_), .S(u5_mult_82_SUMB_40__36_) );
  FA_X1 u5_mult_82_S2_40_35 ( .A(u5_mult_82_ab_40__35_), .B(
        u5_mult_82_CARRYB_39__35_), .CI(u5_mult_82_SUMB_39__36_), .CO(
        u5_mult_82_CARRYB_40__35_), .S(u5_mult_82_SUMB_40__35_) );
  FA_X1 u5_mult_82_S2_40_34 ( .A(u5_mult_82_ab_40__34_), .B(
        u5_mult_82_CARRYB_39__34_), .CI(u5_mult_82_SUMB_39__35_), .CO(
        u5_mult_82_CARRYB_40__34_), .S(u5_mult_82_SUMB_40__34_) );
  FA_X1 u5_mult_82_S2_40_33 ( .A(u5_mult_82_ab_40__33_), .B(
        u5_mult_82_CARRYB_39__33_), .CI(u5_mult_82_SUMB_39__34_), .CO(
        u5_mult_82_CARRYB_40__33_), .S(u5_mult_82_SUMB_40__33_) );
  FA_X1 u5_mult_82_S2_40_32 ( .A(u5_mult_82_ab_40__32_), .B(
        u5_mult_82_CARRYB_39__32_), .CI(u5_mult_82_SUMB_39__33_), .CO(
        u5_mult_82_CARRYB_40__32_), .S(u5_mult_82_SUMB_40__32_) );
  FA_X1 u5_mult_82_S2_40_31 ( .A(u5_mult_82_ab_40__31_), .B(
        u5_mult_82_CARRYB_39__31_), .CI(u5_mult_82_SUMB_39__32_), .CO(
        u5_mult_82_CARRYB_40__31_), .S(u5_mult_82_SUMB_40__31_) );
  FA_X1 u5_mult_82_S2_40_30 ( .A(u5_mult_82_ab_40__30_), .B(
        u5_mult_82_CARRYB_39__30_), .CI(u5_mult_82_SUMB_39__31_), .CO(
        u5_mult_82_CARRYB_40__30_), .S(u5_mult_82_SUMB_40__30_) );
  FA_X1 u5_mult_82_S2_40_29 ( .A(u5_mult_82_ab_40__29_), .B(
        u5_mult_82_CARRYB_39__29_), .CI(u5_mult_82_SUMB_39__30_), .CO(
        u5_mult_82_CARRYB_40__29_), .S(u5_mult_82_SUMB_40__29_) );
  FA_X1 u5_mult_82_S2_40_28 ( .A(u5_mult_82_ab_40__28_), .B(
        u5_mult_82_CARRYB_39__28_), .CI(u5_mult_82_SUMB_39__29_), .CO(
        u5_mult_82_CARRYB_40__28_), .S(u5_mult_82_SUMB_40__28_) );
  FA_X1 u5_mult_82_S2_40_27 ( .A(u5_mult_82_ab_40__27_), .B(
        u5_mult_82_CARRYB_39__27_), .CI(u5_mult_82_SUMB_39__28_), .CO(
        u5_mult_82_CARRYB_40__27_), .S(u5_mult_82_SUMB_40__27_) );
  FA_X1 u5_mult_82_S2_40_26 ( .A(u5_mult_82_ab_40__26_), .B(
        u5_mult_82_CARRYB_39__26_), .CI(u5_mult_82_SUMB_39__27_), .CO(
        u5_mult_82_CARRYB_40__26_), .S(u5_mult_82_SUMB_40__26_) );
  FA_X1 u5_mult_82_S2_40_25 ( .A(u5_mult_82_ab_40__25_), .B(
        u5_mult_82_CARRYB_39__25_), .CI(u5_mult_82_SUMB_39__26_), .CO(
        u5_mult_82_CARRYB_40__25_), .S(u5_mult_82_SUMB_40__25_) );
  FA_X1 u5_mult_82_S2_40_24 ( .A(u5_mult_82_ab_40__24_), .B(
        u5_mult_82_CARRYB_39__24_), .CI(u5_mult_82_SUMB_39__25_), .CO(
        u5_mult_82_CARRYB_40__24_), .S(u5_mult_82_SUMB_40__24_) );
  FA_X1 u5_mult_82_S2_40_23 ( .A(u5_mult_82_ab_40__23_), .B(
        u5_mult_82_CARRYB_39__23_), .CI(u5_mult_82_SUMB_39__24_), .CO(
        u5_mult_82_CARRYB_40__23_), .S(u5_mult_82_SUMB_40__23_) );
  FA_X1 u5_mult_82_S2_40_22 ( .A(u5_mult_82_ab_40__22_), .B(
        u5_mult_82_CARRYB_39__22_), .CI(u5_mult_82_SUMB_39__23_), .CO(
        u5_mult_82_CARRYB_40__22_), .S(u5_mult_82_SUMB_40__22_) );
  FA_X1 u5_mult_82_S2_40_21 ( .A(u5_mult_82_ab_40__21_), .B(
        u5_mult_82_CARRYB_39__21_), .CI(u5_mult_82_SUMB_39__22_), .CO(
        u5_mult_82_CARRYB_40__21_), .S(u5_mult_82_SUMB_40__21_) );
  FA_X1 u5_mult_82_S2_40_20 ( .A(u5_mult_82_ab_40__20_), .B(
        u5_mult_82_CARRYB_39__20_), .CI(u5_mult_82_SUMB_39__21_), .CO(
        u5_mult_82_CARRYB_40__20_), .S(u5_mult_82_SUMB_40__20_) );
  FA_X1 u5_mult_82_S2_40_19 ( .A(u5_mult_82_ab_40__19_), .B(
        u5_mult_82_CARRYB_39__19_), .CI(u5_mult_82_SUMB_39__20_), .CO(
        u5_mult_82_CARRYB_40__19_), .S(u5_mult_82_SUMB_40__19_) );
  FA_X1 u5_mult_82_S2_40_18 ( .A(u5_mult_82_ab_40__18_), .B(
        u5_mult_82_CARRYB_39__18_), .CI(u5_mult_82_SUMB_39__19_), .CO(
        u5_mult_82_CARRYB_40__18_), .S(u5_mult_82_SUMB_40__18_) );
  FA_X1 u5_mult_82_S2_40_17 ( .A(u5_mult_82_ab_40__17_), .B(
        u5_mult_82_CARRYB_39__17_), .CI(u5_mult_82_SUMB_39__18_), .CO(
        u5_mult_82_CARRYB_40__17_), .S(u5_mult_82_SUMB_40__17_) );
  FA_X1 u5_mult_82_S2_40_16 ( .A(u5_mult_82_ab_40__16_), .B(
        u5_mult_82_CARRYB_39__16_), .CI(u5_mult_82_SUMB_39__17_), .CO(
        u5_mult_82_CARRYB_40__16_), .S(u5_mult_82_SUMB_40__16_) );
  FA_X1 u5_mult_82_S2_40_15 ( .A(u5_mult_82_ab_40__15_), .B(
        u5_mult_82_CARRYB_39__15_), .CI(u5_mult_82_SUMB_39__16_), .CO(
        u5_mult_82_CARRYB_40__15_), .S(u5_mult_82_SUMB_40__15_) );
  FA_X1 u5_mult_82_S2_40_14 ( .A(u5_mult_82_ab_40__14_), .B(
        u5_mult_82_CARRYB_39__14_), .CI(u5_mult_82_SUMB_39__15_), .CO(
        u5_mult_82_CARRYB_40__14_), .S(u5_mult_82_SUMB_40__14_) );
  FA_X1 u5_mult_82_S2_40_13 ( .A(u5_mult_82_ab_40__13_), .B(
        u5_mult_82_CARRYB_39__13_), .CI(u5_mult_82_SUMB_39__14_), .CO(
        u5_mult_82_CARRYB_40__13_), .S(u5_mult_82_SUMB_40__13_) );
  FA_X1 u5_mult_82_S2_40_12 ( .A(u5_mult_82_ab_40__12_), .B(
        u5_mult_82_CARRYB_39__12_), .CI(u5_mult_82_SUMB_39__13_), .CO(
        u5_mult_82_CARRYB_40__12_), .S(u5_mult_82_SUMB_40__12_) );
  FA_X1 u5_mult_82_S2_40_11 ( .A(u5_mult_82_ab_40__11_), .B(
        u5_mult_82_CARRYB_39__11_), .CI(u5_mult_82_SUMB_39__12_), .CO(
        u5_mult_82_CARRYB_40__11_), .S(u5_mult_82_SUMB_40__11_) );
  FA_X1 u5_mult_82_S2_40_10 ( .A(u5_mult_82_ab_40__10_), .B(
        u5_mult_82_CARRYB_39__10_), .CI(u5_mult_82_SUMB_39__11_), .CO(
        u5_mult_82_CARRYB_40__10_), .S(u5_mult_82_SUMB_40__10_) );
  FA_X1 u5_mult_82_S2_40_9 ( .A(u5_mult_82_ab_40__9_), .B(
        u5_mult_82_CARRYB_39__9_), .CI(u5_mult_82_SUMB_39__10_), .CO(
        u5_mult_82_CARRYB_40__9_), .S(u5_mult_82_SUMB_40__9_) );
  FA_X1 u5_mult_82_S2_40_8 ( .A(u5_mult_82_ab_40__8_), .B(
        u5_mult_82_CARRYB_39__8_), .CI(u5_mult_82_SUMB_39__9_), .CO(
        u5_mult_82_CARRYB_40__8_), .S(u5_mult_82_SUMB_40__8_) );
  FA_X1 u5_mult_82_S2_40_7 ( .A(u5_mult_82_ab_40__7_), .B(
        u5_mult_82_CARRYB_39__7_), .CI(u5_mult_82_SUMB_39__8_), .CO(
        u5_mult_82_CARRYB_40__7_), .S(u5_mult_82_SUMB_40__7_) );
  FA_X1 u5_mult_82_S2_40_6 ( .A(u5_mult_82_ab_40__6_), .B(
        u5_mult_82_CARRYB_39__6_), .CI(u5_mult_82_SUMB_39__7_), .CO(
        u5_mult_82_CARRYB_40__6_), .S(u5_mult_82_SUMB_40__6_) );
  FA_X1 u5_mult_82_S2_40_5 ( .A(u5_mult_82_ab_40__5_), .B(
        u5_mult_82_CARRYB_39__5_), .CI(u5_mult_82_SUMB_39__6_), .CO(
        u5_mult_82_CARRYB_40__5_), .S(u5_mult_82_SUMB_40__5_) );
  FA_X1 u5_mult_82_S2_40_4 ( .A(u5_mult_82_ab_40__4_), .B(
        u5_mult_82_CARRYB_39__4_), .CI(u5_mult_82_SUMB_39__5_), .CO(
        u5_mult_82_CARRYB_40__4_), .S(u5_mult_82_SUMB_40__4_) );
  FA_X1 u5_mult_82_S2_40_3 ( .A(u5_mult_82_ab_40__3_), .B(
        u5_mult_82_CARRYB_39__3_), .CI(u5_mult_82_SUMB_39__4_), .CO(
        u5_mult_82_CARRYB_40__3_), .S(u5_mult_82_SUMB_40__3_) );
  FA_X1 u5_mult_82_S2_40_2 ( .A(u5_mult_82_ab_40__2_), .B(
        u5_mult_82_CARRYB_39__2_), .CI(u5_mult_82_SUMB_39__3_), .CO(
        u5_mult_82_CARRYB_40__2_), .S(u5_mult_82_SUMB_40__2_) );
  FA_X1 u5_mult_82_S2_40_1 ( .A(u5_mult_82_ab_40__1_), .B(
        u5_mult_82_CARRYB_39__1_), .CI(u5_mult_82_SUMB_39__2_), .CO(
        u5_mult_82_CARRYB_40__1_), .S(u5_mult_82_SUMB_40__1_) );
  FA_X1 u5_mult_82_S1_40_0 ( .A(u5_mult_82_ab_40__0_), .B(
        u5_mult_82_CARRYB_39__0_), .CI(u5_mult_82_SUMB_39__1_), .CO(
        u5_mult_82_CARRYB_40__0_), .S(u5_N40) );
  FA_X1 u5_mult_82_S3_41_51 ( .A(u5_mult_82_ab_41__51_), .B(
        u5_mult_82_CARRYB_40__51_), .CI(u5_mult_82_ab_40__52_), .CO(
        u5_mult_82_CARRYB_41__51_), .S(u5_mult_82_SUMB_41__51_) );
  FA_X1 u5_mult_82_S2_41_50 ( .A(u5_mult_82_ab_41__50_), .B(
        u5_mult_82_CARRYB_40__50_), .CI(u5_mult_82_SUMB_40__51_), .CO(
        u5_mult_82_CARRYB_41__50_), .S(u5_mult_82_SUMB_41__50_) );
  FA_X1 u5_mult_82_S2_41_49 ( .A(u5_mult_82_ab_41__49_), .B(
        u5_mult_82_CARRYB_40__49_), .CI(u5_mult_82_SUMB_40__50_), .CO(
        u5_mult_82_CARRYB_41__49_), .S(u5_mult_82_SUMB_41__49_) );
  FA_X1 u5_mult_82_S2_41_48 ( .A(u5_mult_82_ab_41__48_), .B(
        u5_mult_82_CARRYB_40__48_), .CI(u5_mult_82_SUMB_40__49_), .CO(
        u5_mult_82_CARRYB_41__48_), .S(u5_mult_82_SUMB_41__48_) );
  FA_X1 u5_mult_82_S2_41_47 ( .A(u5_mult_82_ab_41__47_), .B(
        u5_mult_82_CARRYB_40__47_), .CI(u5_mult_82_SUMB_40__48_), .CO(
        u5_mult_82_CARRYB_41__47_), .S(u5_mult_82_SUMB_41__47_) );
  FA_X1 u5_mult_82_S2_41_46 ( .A(u5_mult_82_ab_41__46_), .B(
        u5_mult_82_CARRYB_40__46_), .CI(u5_mult_82_SUMB_40__47_), .CO(
        u5_mult_82_CARRYB_41__46_), .S(u5_mult_82_SUMB_41__46_) );
  FA_X1 u5_mult_82_S2_41_45 ( .A(u5_mult_82_ab_41__45_), .B(
        u5_mult_82_CARRYB_40__45_), .CI(u5_mult_82_SUMB_40__46_), .CO(
        u5_mult_82_CARRYB_41__45_), .S(u5_mult_82_SUMB_41__45_) );
  FA_X1 u5_mult_82_S2_41_44 ( .A(u5_mult_82_ab_41__44_), .B(
        u5_mult_82_CARRYB_40__44_), .CI(u5_mult_82_SUMB_40__45_), .CO(
        u5_mult_82_CARRYB_41__44_), .S(u5_mult_82_SUMB_41__44_) );
  FA_X1 u5_mult_82_S2_41_43 ( .A(u5_mult_82_ab_41__43_), .B(
        u5_mult_82_CARRYB_40__43_), .CI(u5_mult_82_SUMB_40__44_), .CO(
        u5_mult_82_CARRYB_41__43_), .S(u5_mult_82_SUMB_41__43_) );
  FA_X1 u5_mult_82_S2_41_42 ( .A(u5_mult_82_ab_41__42_), .B(
        u5_mult_82_CARRYB_40__42_), .CI(u5_mult_82_SUMB_40__43_), .CO(
        u5_mult_82_CARRYB_41__42_), .S(u5_mult_82_SUMB_41__42_) );
  FA_X1 u5_mult_82_S2_41_41 ( .A(u5_mult_82_ab_41__41_), .B(
        u5_mult_82_CARRYB_40__41_), .CI(u5_mult_82_SUMB_40__42_), .CO(
        u5_mult_82_CARRYB_41__41_), .S(u5_mult_82_SUMB_41__41_) );
  FA_X1 u5_mult_82_S2_41_40 ( .A(u5_mult_82_ab_41__40_), .B(
        u5_mult_82_CARRYB_40__40_), .CI(u5_mult_82_SUMB_40__41_), .CO(
        u5_mult_82_CARRYB_41__40_), .S(u5_mult_82_SUMB_41__40_) );
  FA_X1 u5_mult_82_S2_41_39 ( .A(u5_mult_82_ab_41__39_), .B(
        u5_mult_82_CARRYB_40__39_), .CI(u5_mult_82_SUMB_40__40_), .CO(
        u5_mult_82_CARRYB_41__39_), .S(u5_mult_82_SUMB_41__39_) );
  FA_X1 u5_mult_82_S2_41_38 ( .A(u5_mult_82_ab_41__38_), .B(
        u5_mult_82_CARRYB_40__38_), .CI(u5_mult_82_SUMB_40__39_), .CO(
        u5_mult_82_CARRYB_41__38_), .S(u5_mult_82_SUMB_41__38_) );
  FA_X1 u5_mult_82_S2_41_37 ( .A(u5_mult_82_ab_41__37_), .B(
        u5_mult_82_CARRYB_40__37_), .CI(u5_mult_82_SUMB_40__38_), .CO(
        u5_mult_82_CARRYB_41__37_), .S(u5_mult_82_SUMB_41__37_) );
  FA_X1 u5_mult_82_S2_41_36 ( .A(u5_mult_82_ab_41__36_), .B(
        u5_mult_82_CARRYB_40__36_), .CI(u5_mult_82_SUMB_40__37_), .CO(
        u5_mult_82_CARRYB_41__36_), .S(u5_mult_82_SUMB_41__36_) );
  FA_X1 u5_mult_82_S2_41_35 ( .A(u5_mult_82_ab_41__35_), .B(
        u5_mult_82_CARRYB_40__35_), .CI(u5_mult_82_SUMB_40__36_), .CO(
        u5_mult_82_CARRYB_41__35_), .S(u5_mult_82_SUMB_41__35_) );
  FA_X1 u5_mult_82_S2_41_34 ( .A(u5_mult_82_ab_41__34_), .B(
        u5_mult_82_CARRYB_40__34_), .CI(u5_mult_82_SUMB_40__35_), .CO(
        u5_mult_82_CARRYB_41__34_), .S(u5_mult_82_SUMB_41__34_) );
  FA_X1 u5_mult_82_S2_41_33 ( .A(u5_mult_82_ab_41__33_), .B(
        u5_mult_82_CARRYB_40__33_), .CI(u5_mult_82_SUMB_40__34_), .CO(
        u5_mult_82_CARRYB_41__33_), .S(u5_mult_82_SUMB_41__33_) );
  FA_X1 u5_mult_82_S2_41_32 ( .A(u5_mult_82_ab_41__32_), .B(
        u5_mult_82_CARRYB_40__32_), .CI(u5_mult_82_SUMB_40__33_), .CO(
        u5_mult_82_CARRYB_41__32_), .S(u5_mult_82_SUMB_41__32_) );
  FA_X1 u5_mult_82_S2_41_31 ( .A(u5_mult_82_ab_41__31_), .B(
        u5_mult_82_CARRYB_40__31_), .CI(u5_mult_82_SUMB_40__32_), .CO(
        u5_mult_82_CARRYB_41__31_), .S(u5_mult_82_SUMB_41__31_) );
  FA_X1 u5_mult_82_S2_41_30 ( .A(u5_mult_82_ab_41__30_), .B(
        u5_mult_82_CARRYB_40__30_), .CI(u5_mult_82_SUMB_40__31_), .CO(
        u5_mult_82_CARRYB_41__30_), .S(u5_mult_82_SUMB_41__30_) );
  FA_X1 u5_mult_82_S2_41_29 ( .A(u5_mult_82_ab_41__29_), .B(
        u5_mult_82_CARRYB_40__29_), .CI(u5_mult_82_SUMB_40__30_), .CO(
        u5_mult_82_CARRYB_41__29_), .S(u5_mult_82_SUMB_41__29_) );
  FA_X1 u5_mult_82_S2_41_28 ( .A(u5_mult_82_ab_41__28_), .B(
        u5_mult_82_CARRYB_40__28_), .CI(u5_mult_82_SUMB_40__29_), .CO(
        u5_mult_82_CARRYB_41__28_), .S(u5_mult_82_SUMB_41__28_) );
  FA_X1 u5_mult_82_S2_41_27 ( .A(u5_mult_82_ab_41__27_), .B(
        u5_mult_82_CARRYB_40__27_), .CI(u5_mult_82_SUMB_40__28_), .CO(
        u5_mult_82_CARRYB_41__27_), .S(u5_mult_82_SUMB_41__27_) );
  FA_X1 u5_mult_82_S2_41_26 ( .A(u5_mult_82_ab_41__26_), .B(
        u5_mult_82_CARRYB_40__26_), .CI(u5_mult_82_SUMB_40__27_), .CO(
        u5_mult_82_CARRYB_41__26_), .S(u5_mult_82_SUMB_41__26_) );
  FA_X1 u5_mult_82_S2_41_25 ( .A(u5_mult_82_ab_41__25_), .B(
        u5_mult_82_CARRYB_40__25_), .CI(u5_mult_82_SUMB_40__26_), .CO(
        u5_mult_82_CARRYB_41__25_), .S(u5_mult_82_SUMB_41__25_) );
  FA_X1 u5_mult_82_S2_41_24 ( .A(u5_mult_82_ab_41__24_), .B(
        u5_mult_82_CARRYB_40__24_), .CI(u5_mult_82_SUMB_40__25_), .CO(
        u5_mult_82_CARRYB_41__24_), .S(u5_mult_82_SUMB_41__24_) );
  FA_X1 u5_mult_82_S2_41_23 ( .A(u5_mult_82_ab_41__23_), .B(
        u5_mult_82_CARRYB_40__23_), .CI(u5_mult_82_SUMB_40__24_), .CO(
        u5_mult_82_CARRYB_41__23_), .S(u5_mult_82_SUMB_41__23_) );
  FA_X1 u5_mult_82_S2_41_22 ( .A(u5_mult_82_ab_41__22_), .B(
        u5_mult_82_CARRYB_40__22_), .CI(u5_mult_82_SUMB_40__23_), .CO(
        u5_mult_82_CARRYB_41__22_), .S(u5_mult_82_SUMB_41__22_) );
  FA_X1 u5_mult_82_S2_41_21 ( .A(u5_mult_82_ab_41__21_), .B(
        u5_mult_82_CARRYB_40__21_), .CI(u5_mult_82_SUMB_40__22_), .CO(
        u5_mult_82_CARRYB_41__21_), .S(u5_mult_82_SUMB_41__21_) );
  FA_X1 u5_mult_82_S2_41_20 ( .A(u5_mult_82_ab_41__20_), .B(
        u5_mult_82_CARRYB_40__20_), .CI(u5_mult_82_SUMB_40__21_), .CO(
        u5_mult_82_CARRYB_41__20_), .S(u5_mult_82_SUMB_41__20_) );
  FA_X1 u5_mult_82_S2_41_19 ( .A(u5_mult_82_ab_41__19_), .B(
        u5_mult_82_CARRYB_40__19_), .CI(u5_mult_82_SUMB_40__20_), .CO(
        u5_mult_82_CARRYB_41__19_), .S(u5_mult_82_SUMB_41__19_) );
  FA_X1 u5_mult_82_S2_41_18 ( .A(u5_mult_82_ab_41__18_), .B(
        u5_mult_82_CARRYB_40__18_), .CI(u5_mult_82_SUMB_40__19_), .CO(
        u5_mult_82_CARRYB_41__18_), .S(u5_mult_82_SUMB_41__18_) );
  FA_X1 u5_mult_82_S2_41_17 ( .A(u5_mult_82_ab_41__17_), .B(
        u5_mult_82_CARRYB_40__17_), .CI(u5_mult_82_SUMB_40__18_), .CO(
        u5_mult_82_CARRYB_41__17_), .S(u5_mult_82_SUMB_41__17_) );
  FA_X1 u5_mult_82_S2_41_16 ( .A(u5_mult_82_ab_41__16_), .B(
        u5_mult_82_CARRYB_40__16_), .CI(u5_mult_82_SUMB_40__17_), .CO(
        u5_mult_82_CARRYB_41__16_), .S(u5_mult_82_SUMB_41__16_) );
  FA_X1 u5_mult_82_S2_41_15 ( .A(u5_mult_82_ab_41__15_), .B(
        u5_mult_82_CARRYB_40__15_), .CI(u5_mult_82_SUMB_40__16_), .CO(
        u5_mult_82_CARRYB_41__15_), .S(u5_mult_82_SUMB_41__15_) );
  FA_X1 u5_mult_82_S2_41_14 ( .A(u5_mult_82_ab_41__14_), .B(
        u5_mult_82_CARRYB_40__14_), .CI(u5_mult_82_SUMB_40__15_), .CO(
        u5_mult_82_CARRYB_41__14_), .S(u5_mult_82_SUMB_41__14_) );
  FA_X1 u5_mult_82_S2_41_13 ( .A(u5_mult_82_ab_41__13_), .B(
        u5_mult_82_CARRYB_40__13_), .CI(u5_mult_82_SUMB_40__14_), .CO(
        u5_mult_82_CARRYB_41__13_), .S(u5_mult_82_SUMB_41__13_) );
  FA_X1 u5_mult_82_S2_41_12 ( .A(u5_mult_82_ab_41__12_), .B(
        u5_mult_82_CARRYB_40__12_), .CI(u5_mult_82_SUMB_40__13_), .CO(
        u5_mult_82_CARRYB_41__12_), .S(u5_mult_82_SUMB_41__12_) );
  FA_X1 u5_mult_82_S2_41_11 ( .A(u5_mult_82_ab_41__11_), .B(
        u5_mult_82_CARRYB_40__11_), .CI(u5_mult_82_SUMB_40__12_), .CO(
        u5_mult_82_CARRYB_41__11_), .S(u5_mult_82_SUMB_41__11_) );
  FA_X1 u5_mult_82_S2_41_10 ( .A(u5_mult_82_ab_41__10_), .B(
        u5_mult_82_CARRYB_40__10_), .CI(u5_mult_82_SUMB_40__11_), .CO(
        u5_mult_82_CARRYB_41__10_), .S(u5_mult_82_SUMB_41__10_) );
  FA_X1 u5_mult_82_S2_41_9 ( .A(u5_mult_82_ab_41__9_), .B(
        u5_mult_82_CARRYB_40__9_), .CI(u5_mult_82_SUMB_40__10_), .CO(
        u5_mult_82_CARRYB_41__9_), .S(u5_mult_82_SUMB_41__9_) );
  FA_X1 u5_mult_82_S2_41_8 ( .A(u5_mult_82_ab_41__8_), .B(
        u5_mult_82_CARRYB_40__8_), .CI(u5_mult_82_SUMB_40__9_), .CO(
        u5_mult_82_CARRYB_41__8_), .S(u5_mult_82_SUMB_41__8_) );
  FA_X1 u5_mult_82_S2_41_7 ( .A(u5_mult_82_ab_41__7_), .B(
        u5_mult_82_CARRYB_40__7_), .CI(u5_mult_82_SUMB_40__8_), .CO(
        u5_mult_82_CARRYB_41__7_), .S(u5_mult_82_SUMB_41__7_) );
  FA_X1 u5_mult_82_S2_41_6 ( .A(u5_mult_82_ab_41__6_), .B(
        u5_mult_82_CARRYB_40__6_), .CI(u5_mult_82_SUMB_40__7_), .CO(
        u5_mult_82_CARRYB_41__6_), .S(u5_mult_82_SUMB_41__6_) );
  FA_X1 u5_mult_82_S2_41_5 ( .A(u5_mult_82_ab_41__5_), .B(
        u5_mult_82_CARRYB_40__5_), .CI(u5_mult_82_SUMB_40__6_), .CO(
        u5_mult_82_CARRYB_41__5_), .S(u5_mult_82_SUMB_41__5_) );
  FA_X1 u5_mult_82_S2_41_4 ( .A(u5_mult_82_ab_41__4_), .B(
        u5_mult_82_CARRYB_40__4_), .CI(u5_mult_82_SUMB_40__5_), .CO(
        u5_mult_82_CARRYB_41__4_), .S(u5_mult_82_SUMB_41__4_) );
  FA_X1 u5_mult_82_S2_41_3 ( .A(u5_mult_82_ab_41__3_), .B(
        u5_mult_82_CARRYB_40__3_), .CI(u5_mult_82_SUMB_40__4_), .CO(
        u5_mult_82_CARRYB_41__3_), .S(u5_mult_82_SUMB_41__3_) );
  FA_X1 u5_mult_82_S2_41_2 ( .A(u5_mult_82_ab_41__2_), .B(
        u5_mult_82_CARRYB_40__2_), .CI(u5_mult_82_SUMB_40__3_), .CO(
        u5_mult_82_CARRYB_41__2_), .S(u5_mult_82_SUMB_41__2_) );
  FA_X1 u5_mult_82_S2_41_1 ( .A(u5_mult_82_ab_41__1_), .B(
        u5_mult_82_CARRYB_40__1_), .CI(u5_mult_82_SUMB_40__2_), .CO(
        u5_mult_82_CARRYB_41__1_), .S(u5_mult_82_SUMB_41__1_) );
  FA_X1 u5_mult_82_S1_41_0 ( .A(u5_mult_82_ab_41__0_), .B(
        u5_mult_82_CARRYB_40__0_), .CI(u5_mult_82_SUMB_40__1_), .CO(
        u5_mult_82_CARRYB_41__0_), .S(u5_N41) );
  FA_X1 u5_mult_82_S3_42_51 ( .A(u5_mult_82_ab_42__51_), .B(
        u5_mult_82_CARRYB_41__51_), .CI(u5_mult_82_ab_41__52_), .CO(
        u5_mult_82_CARRYB_42__51_), .S(u5_mult_82_SUMB_42__51_) );
  FA_X1 u5_mult_82_S2_42_50 ( .A(u5_mult_82_ab_42__50_), .B(
        u5_mult_82_CARRYB_41__50_), .CI(u5_mult_82_SUMB_41__51_), .CO(
        u5_mult_82_CARRYB_42__50_), .S(u5_mult_82_SUMB_42__50_) );
  FA_X1 u5_mult_82_S2_42_49 ( .A(u5_mult_82_ab_42__49_), .B(
        u5_mult_82_CARRYB_41__49_), .CI(u5_mult_82_SUMB_41__50_), .CO(
        u5_mult_82_CARRYB_42__49_), .S(u5_mult_82_SUMB_42__49_) );
  FA_X1 u5_mult_82_S2_42_48 ( .A(u5_mult_82_ab_42__48_), .B(
        u5_mult_82_CARRYB_41__48_), .CI(u5_mult_82_SUMB_41__49_), .CO(
        u5_mult_82_CARRYB_42__48_), .S(u5_mult_82_SUMB_42__48_) );
  FA_X1 u5_mult_82_S2_42_47 ( .A(u5_mult_82_ab_42__47_), .B(
        u5_mult_82_CARRYB_41__47_), .CI(u5_mult_82_SUMB_41__48_), .CO(
        u5_mult_82_CARRYB_42__47_), .S(u5_mult_82_SUMB_42__47_) );
  FA_X1 u5_mult_82_S2_42_46 ( .A(u5_mult_82_ab_42__46_), .B(
        u5_mult_82_CARRYB_41__46_), .CI(u5_mult_82_SUMB_41__47_), .CO(
        u5_mult_82_CARRYB_42__46_), .S(u5_mult_82_SUMB_42__46_) );
  FA_X1 u5_mult_82_S2_42_45 ( .A(u5_mult_82_ab_42__45_), .B(
        u5_mult_82_CARRYB_41__45_), .CI(u5_mult_82_SUMB_41__46_), .CO(
        u5_mult_82_CARRYB_42__45_), .S(u5_mult_82_SUMB_42__45_) );
  FA_X1 u5_mult_82_S2_42_44 ( .A(u5_mult_82_ab_42__44_), .B(
        u5_mult_82_CARRYB_41__44_), .CI(u5_mult_82_SUMB_41__45_), .CO(
        u5_mult_82_CARRYB_42__44_), .S(u5_mult_82_SUMB_42__44_) );
  FA_X1 u5_mult_82_S2_42_43 ( .A(u5_mult_82_ab_42__43_), .B(
        u5_mult_82_CARRYB_41__43_), .CI(u5_mult_82_SUMB_41__44_), .CO(
        u5_mult_82_CARRYB_42__43_), .S(u5_mult_82_SUMB_42__43_) );
  FA_X1 u5_mult_82_S2_42_42 ( .A(u5_mult_82_ab_42__42_), .B(
        u5_mult_82_CARRYB_41__42_), .CI(u5_mult_82_SUMB_41__43_), .CO(
        u5_mult_82_CARRYB_42__42_), .S(u5_mult_82_SUMB_42__42_) );
  FA_X1 u5_mult_82_S2_42_41 ( .A(u5_mult_82_ab_42__41_), .B(
        u5_mult_82_CARRYB_41__41_), .CI(u5_mult_82_SUMB_41__42_), .CO(
        u5_mult_82_CARRYB_42__41_), .S(u5_mult_82_SUMB_42__41_) );
  FA_X1 u5_mult_82_S2_42_40 ( .A(u5_mult_82_ab_42__40_), .B(
        u5_mult_82_CARRYB_41__40_), .CI(u5_mult_82_SUMB_41__41_), .CO(
        u5_mult_82_CARRYB_42__40_), .S(u5_mult_82_SUMB_42__40_) );
  FA_X1 u5_mult_82_S2_42_39 ( .A(u5_mult_82_ab_42__39_), .B(
        u5_mult_82_CARRYB_41__39_), .CI(u5_mult_82_SUMB_41__40_), .CO(
        u5_mult_82_CARRYB_42__39_), .S(u5_mult_82_SUMB_42__39_) );
  FA_X1 u5_mult_82_S2_42_38 ( .A(u5_mult_82_ab_42__38_), .B(
        u5_mult_82_CARRYB_41__38_), .CI(u5_mult_82_SUMB_41__39_), .CO(
        u5_mult_82_CARRYB_42__38_), .S(u5_mult_82_SUMB_42__38_) );
  FA_X1 u5_mult_82_S2_42_37 ( .A(u5_mult_82_ab_42__37_), .B(
        u5_mult_82_CARRYB_41__37_), .CI(u5_mult_82_SUMB_41__38_), .CO(
        u5_mult_82_CARRYB_42__37_), .S(u5_mult_82_SUMB_42__37_) );
  FA_X1 u5_mult_82_S2_42_36 ( .A(u5_mult_82_ab_42__36_), .B(
        u5_mult_82_CARRYB_41__36_), .CI(u5_mult_82_SUMB_41__37_), .CO(
        u5_mult_82_CARRYB_42__36_), .S(u5_mult_82_SUMB_42__36_) );
  FA_X1 u5_mult_82_S2_42_35 ( .A(u5_mult_82_ab_42__35_), .B(
        u5_mult_82_CARRYB_41__35_), .CI(u5_mult_82_SUMB_41__36_), .CO(
        u5_mult_82_CARRYB_42__35_), .S(u5_mult_82_SUMB_42__35_) );
  FA_X1 u5_mult_82_S2_42_34 ( .A(u5_mult_82_ab_42__34_), .B(
        u5_mult_82_CARRYB_41__34_), .CI(u5_mult_82_SUMB_41__35_), .CO(
        u5_mult_82_CARRYB_42__34_), .S(u5_mult_82_SUMB_42__34_) );
  FA_X1 u5_mult_82_S2_42_33 ( .A(u5_mult_82_ab_42__33_), .B(
        u5_mult_82_CARRYB_41__33_), .CI(u5_mult_82_SUMB_41__34_), .CO(
        u5_mult_82_CARRYB_42__33_), .S(u5_mult_82_SUMB_42__33_) );
  FA_X1 u5_mult_82_S2_42_32 ( .A(u5_mult_82_ab_42__32_), .B(
        u5_mult_82_CARRYB_41__32_), .CI(u5_mult_82_SUMB_41__33_), .CO(
        u5_mult_82_CARRYB_42__32_), .S(u5_mult_82_SUMB_42__32_) );
  FA_X1 u5_mult_82_S2_42_31 ( .A(u5_mult_82_ab_42__31_), .B(
        u5_mult_82_CARRYB_41__31_), .CI(u5_mult_82_SUMB_41__32_), .CO(
        u5_mult_82_CARRYB_42__31_), .S(u5_mult_82_SUMB_42__31_) );
  FA_X1 u5_mult_82_S2_42_30 ( .A(u5_mult_82_ab_42__30_), .B(
        u5_mult_82_CARRYB_41__30_), .CI(u5_mult_82_SUMB_41__31_), .CO(
        u5_mult_82_CARRYB_42__30_), .S(u5_mult_82_SUMB_42__30_) );
  FA_X1 u5_mult_82_S2_42_29 ( .A(u5_mult_82_ab_42__29_), .B(
        u5_mult_82_CARRYB_41__29_), .CI(u5_mult_82_SUMB_41__30_), .CO(
        u5_mult_82_CARRYB_42__29_), .S(u5_mult_82_SUMB_42__29_) );
  FA_X1 u5_mult_82_S2_42_28 ( .A(u5_mult_82_ab_42__28_), .B(
        u5_mult_82_CARRYB_41__28_), .CI(u5_mult_82_SUMB_41__29_), .CO(
        u5_mult_82_CARRYB_42__28_), .S(u5_mult_82_SUMB_42__28_) );
  FA_X1 u5_mult_82_S2_42_27 ( .A(u5_mult_82_ab_42__27_), .B(
        u5_mult_82_CARRYB_41__27_), .CI(u5_mult_82_SUMB_41__28_), .CO(
        u5_mult_82_CARRYB_42__27_), .S(u5_mult_82_SUMB_42__27_) );
  FA_X1 u5_mult_82_S2_42_26 ( .A(u5_mult_82_ab_42__26_), .B(
        u5_mult_82_CARRYB_41__26_), .CI(u5_mult_82_SUMB_41__27_), .CO(
        u5_mult_82_CARRYB_42__26_), .S(u5_mult_82_SUMB_42__26_) );
  FA_X1 u5_mult_82_S2_42_25 ( .A(u5_mult_82_ab_42__25_), .B(
        u5_mult_82_CARRYB_41__25_), .CI(u5_mult_82_SUMB_41__26_), .CO(
        u5_mult_82_CARRYB_42__25_), .S(u5_mult_82_SUMB_42__25_) );
  FA_X1 u5_mult_82_S2_42_24 ( .A(u5_mult_82_ab_42__24_), .B(
        u5_mult_82_CARRYB_41__24_), .CI(u5_mult_82_SUMB_41__25_), .CO(
        u5_mult_82_CARRYB_42__24_), .S(u5_mult_82_SUMB_42__24_) );
  FA_X1 u5_mult_82_S2_42_23 ( .A(u5_mult_82_ab_42__23_), .B(
        u5_mult_82_CARRYB_41__23_), .CI(u5_mult_82_SUMB_41__24_), .CO(
        u5_mult_82_CARRYB_42__23_), .S(u5_mult_82_SUMB_42__23_) );
  FA_X1 u5_mult_82_S2_42_22 ( .A(u5_mult_82_ab_42__22_), .B(
        u5_mult_82_CARRYB_41__22_), .CI(u5_mult_82_SUMB_41__23_), .CO(
        u5_mult_82_CARRYB_42__22_), .S(u5_mult_82_SUMB_42__22_) );
  FA_X1 u5_mult_82_S2_42_21 ( .A(u5_mult_82_ab_42__21_), .B(
        u5_mult_82_CARRYB_41__21_), .CI(u5_mult_82_SUMB_41__22_), .CO(
        u5_mult_82_CARRYB_42__21_), .S(u5_mult_82_SUMB_42__21_) );
  FA_X1 u5_mult_82_S2_42_20 ( .A(u5_mult_82_ab_42__20_), .B(
        u5_mult_82_CARRYB_41__20_), .CI(u5_mult_82_SUMB_41__21_), .CO(
        u5_mult_82_CARRYB_42__20_), .S(u5_mult_82_SUMB_42__20_) );
  FA_X1 u5_mult_82_S2_42_19 ( .A(u5_mult_82_ab_42__19_), .B(
        u5_mult_82_CARRYB_41__19_), .CI(u5_mult_82_SUMB_41__20_), .CO(
        u5_mult_82_CARRYB_42__19_), .S(u5_mult_82_SUMB_42__19_) );
  FA_X1 u5_mult_82_S2_42_18 ( .A(u5_mult_82_ab_42__18_), .B(
        u5_mult_82_CARRYB_41__18_), .CI(u5_mult_82_SUMB_41__19_), .CO(
        u5_mult_82_CARRYB_42__18_), .S(u5_mult_82_SUMB_42__18_) );
  FA_X1 u5_mult_82_S2_42_17 ( .A(u5_mult_82_ab_42__17_), .B(
        u5_mult_82_CARRYB_41__17_), .CI(u5_mult_82_SUMB_41__18_), .CO(
        u5_mult_82_CARRYB_42__17_), .S(u5_mult_82_SUMB_42__17_) );
  FA_X1 u5_mult_82_S2_42_16 ( .A(u5_mult_82_ab_42__16_), .B(
        u5_mult_82_CARRYB_41__16_), .CI(u5_mult_82_SUMB_41__17_), .CO(
        u5_mult_82_CARRYB_42__16_), .S(u5_mult_82_SUMB_42__16_) );
  FA_X1 u5_mult_82_S2_42_15 ( .A(u5_mult_82_ab_42__15_), .B(
        u5_mult_82_CARRYB_41__15_), .CI(u5_mult_82_SUMB_41__16_), .CO(
        u5_mult_82_CARRYB_42__15_), .S(u5_mult_82_SUMB_42__15_) );
  FA_X1 u5_mult_82_S2_42_14 ( .A(u5_mult_82_ab_42__14_), .B(
        u5_mult_82_CARRYB_41__14_), .CI(u5_mult_82_SUMB_41__15_), .CO(
        u5_mult_82_CARRYB_42__14_), .S(u5_mult_82_SUMB_42__14_) );
  FA_X1 u5_mult_82_S2_42_13 ( .A(u5_mult_82_ab_42__13_), .B(
        u5_mult_82_CARRYB_41__13_), .CI(u5_mult_82_SUMB_41__14_), .CO(
        u5_mult_82_CARRYB_42__13_), .S(u5_mult_82_SUMB_42__13_) );
  FA_X1 u5_mult_82_S2_42_12 ( .A(u5_mult_82_ab_42__12_), .B(
        u5_mult_82_CARRYB_41__12_), .CI(u5_mult_82_SUMB_41__13_), .CO(
        u5_mult_82_CARRYB_42__12_), .S(u5_mult_82_SUMB_42__12_) );
  FA_X1 u5_mult_82_S2_42_11 ( .A(u5_mult_82_ab_42__11_), .B(
        u5_mult_82_CARRYB_41__11_), .CI(u5_mult_82_SUMB_41__12_), .CO(
        u5_mult_82_CARRYB_42__11_), .S(u5_mult_82_SUMB_42__11_) );
  FA_X1 u5_mult_82_S2_42_10 ( .A(u5_mult_82_ab_42__10_), .B(
        u5_mult_82_CARRYB_41__10_), .CI(u5_mult_82_SUMB_41__11_), .CO(
        u5_mult_82_CARRYB_42__10_), .S(u5_mult_82_SUMB_42__10_) );
  FA_X1 u5_mult_82_S2_42_9 ( .A(u5_mult_82_ab_42__9_), .B(
        u5_mult_82_CARRYB_41__9_), .CI(u5_mult_82_SUMB_41__10_), .CO(
        u5_mult_82_CARRYB_42__9_), .S(u5_mult_82_SUMB_42__9_) );
  FA_X1 u5_mult_82_S2_42_8 ( .A(u5_mult_82_ab_42__8_), .B(
        u5_mult_82_CARRYB_41__8_), .CI(u5_mult_82_SUMB_41__9_), .CO(
        u5_mult_82_CARRYB_42__8_), .S(u5_mult_82_SUMB_42__8_) );
  FA_X1 u5_mult_82_S2_42_7 ( .A(u5_mult_82_ab_42__7_), .B(
        u5_mult_82_CARRYB_41__7_), .CI(u5_mult_82_SUMB_41__8_), .CO(
        u5_mult_82_CARRYB_42__7_), .S(u5_mult_82_SUMB_42__7_) );
  FA_X1 u5_mult_82_S2_42_6 ( .A(u5_mult_82_ab_42__6_), .B(
        u5_mult_82_CARRYB_41__6_), .CI(u5_mult_82_SUMB_41__7_), .CO(
        u5_mult_82_CARRYB_42__6_), .S(u5_mult_82_SUMB_42__6_) );
  FA_X1 u5_mult_82_S2_42_5 ( .A(u5_mult_82_ab_42__5_), .B(
        u5_mult_82_CARRYB_41__5_), .CI(u5_mult_82_SUMB_41__6_), .CO(
        u5_mult_82_CARRYB_42__5_), .S(u5_mult_82_SUMB_42__5_) );
  FA_X1 u5_mult_82_S2_42_4 ( .A(u5_mult_82_ab_42__4_), .B(
        u5_mult_82_CARRYB_41__4_), .CI(u5_mult_82_SUMB_41__5_), .CO(
        u5_mult_82_CARRYB_42__4_), .S(u5_mult_82_SUMB_42__4_) );
  FA_X1 u5_mult_82_S2_42_3 ( .A(u5_mult_82_ab_42__3_), .B(
        u5_mult_82_CARRYB_41__3_), .CI(u5_mult_82_SUMB_41__4_), .CO(
        u5_mult_82_CARRYB_42__3_), .S(u5_mult_82_SUMB_42__3_) );
  FA_X1 u5_mult_82_S2_42_2 ( .A(u5_mult_82_ab_42__2_), .B(
        u5_mult_82_CARRYB_41__2_), .CI(u5_mult_82_SUMB_41__3_), .CO(
        u5_mult_82_CARRYB_42__2_), .S(u5_mult_82_SUMB_42__2_) );
  FA_X1 u5_mult_82_S2_42_1 ( .A(u5_mult_82_ab_42__1_), .B(
        u5_mult_82_CARRYB_41__1_), .CI(u5_mult_82_SUMB_41__2_), .CO(
        u5_mult_82_CARRYB_42__1_), .S(u5_mult_82_SUMB_42__1_) );
  FA_X1 u5_mult_82_S1_42_0 ( .A(u5_mult_82_ab_42__0_), .B(
        u5_mult_82_CARRYB_41__0_), .CI(u5_mult_82_SUMB_41__1_), .CO(
        u5_mult_82_CARRYB_42__0_), .S(u5_N42) );
  FA_X1 u5_mult_82_S3_43_51 ( .A(u5_mult_82_ab_43__51_), .B(
        u5_mult_82_CARRYB_42__51_), .CI(u5_mult_82_ab_42__52_), .CO(
        u5_mult_82_CARRYB_43__51_), .S(u5_mult_82_SUMB_43__51_) );
  FA_X1 u5_mult_82_S2_43_50 ( .A(u5_mult_82_ab_43__50_), .B(
        u5_mult_82_CARRYB_42__50_), .CI(u5_mult_82_SUMB_42__51_), .CO(
        u5_mult_82_CARRYB_43__50_), .S(u5_mult_82_SUMB_43__50_) );
  FA_X1 u5_mult_82_S2_43_49 ( .A(u5_mult_82_ab_43__49_), .B(
        u5_mult_82_CARRYB_42__49_), .CI(u5_mult_82_SUMB_42__50_), .CO(
        u5_mult_82_CARRYB_43__49_), .S(u5_mult_82_SUMB_43__49_) );
  FA_X1 u5_mult_82_S2_43_48 ( .A(u5_mult_82_ab_43__48_), .B(
        u5_mult_82_CARRYB_42__48_), .CI(u5_mult_82_SUMB_42__49_), .CO(
        u5_mult_82_CARRYB_43__48_), .S(u5_mult_82_SUMB_43__48_) );
  FA_X1 u5_mult_82_S2_43_47 ( .A(u5_mult_82_ab_43__47_), .B(
        u5_mult_82_CARRYB_42__47_), .CI(u5_mult_82_SUMB_42__48_), .CO(
        u5_mult_82_CARRYB_43__47_), .S(u5_mult_82_SUMB_43__47_) );
  FA_X1 u5_mult_82_S2_43_46 ( .A(u5_mult_82_ab_43__46_), .B(
        u5_mult_82_CARRYB_42__46_), .CI(u5_mult_82_SUMB_42__47_), .CO(
        u5_mult_82_CARRYB_43__46_), .S(u5_mult_82_SUMB_43__46_) );
  FA_X1 u5_mult_82_S2_43_45 ( .A(u5_mult_82_ab_43__45_), .B(
        u5_mult_82_CARRYB_42__45_), .CI(u5_mult_82_SUMB_42__46_), .CO(
        u5_mult_82_CARRYB_43__45_), .S(u5_mult_82_SUMB_43__45_) );
  FA_X1 u5_mult_82_S2_43_44 ( .A(u5_mult_82_ab_43__44_), .B(
        u5_mult_82_CARRYB_42__44_), .CI(u5_mult_82_SUMB_42__45_), .CO(
        u5_mult_82_CARRYB_43__44_), .S(u5_mult_82_SUMB_43__44_) );
  FA_X1 u5_mult_82_S2_43_43 ( .A(u5_mult_82_ab_43__43_), .B(
        u5_mult_82_CARRYB_42__43_), .CI(u5_mult_82_SUMB_42__44_), .CO(
        u5_mult_82_CARRYB_43__43_), .S(u5_mult_82_SUMB_43__43_) );
  FA_X1 u5_mult_82_S2_43_42 ( .A(u5_mult_82_ab_43__42_), .B(
        u5_mult_82_CARRYB_42__42_), .CI(u5_mult_82_SUMB_42__43_), .CO(
        u5_mult_82_CARRYB_43__42_), .S(u5_mult_82_SUMB_43__42_) );
  FA_X1 u5_mult_82_S2_43_41 ( .A(u5_mult_82_ab_43__41_), .B(
        u5_mult_82_CARRYB_42__41_), .CI(u5_mult_82_SUMB_42__42_), .CO(
        u5_mult_82_CARRYB_43__41_), .S(u5_mult_82_SUMB_43__41_) );
  FA_X1 u5_mult_82_S2_43_40 ( .A(u5_mult_82_ab_43__40_), .B(
        u5_mult_82_CARRYB_42__40_), .CI(u5_mult_82_SUMB_42__41_), .CO(
        u5_mult_82_CARRYB_43__40_), .S(u5_mult_82_SUMB_43__40_) );
  FA_X1 u5_mult_82_S2_43_39 ( .A(u5_mult_82_ab_43__39_), .B(
        u5_mult_82_CARRYB_42__39_), .CI(u5_mult_82_SUMB_42__40_), .CO(
        u5_mult_82_CARRYB_43__39_), .S(u5_mult_82_SUMB_43__39_) );
  FA_X1 u5_mult_82_S2_43_38 ( .A(u5_mult_82_ab_43__38_), .B(
        u5_mult_82_CARRYB_42__38_), .CI(u5_mult_82_SUMB_42__39_), .CO(
        u5_mult_82_CARRYB_43__38_), .S(u5_mult_82_SUMB_43__38_) );
  FA_X1 u5_mult_82_S2_43_37 ( .A(u5_mult_82_ab_43__37_), .B(
        u5_mult_82_CARRYB_42__37_), .CI(u5_mult_82_SUMB_42__38_), .CO(
        u5_mult_82_CARRYB_43__37_), .S(u5_mult_82_SUMB_43__37_) );
  FA_X1 u5_mult_82_S2_43_36 ( .A(u5_mult_82_ab_43__36_), .B(
        u5_mult_82_CARRYB_42__36_), .CI(u5_mult_82_SUMB_42__37_), .CO(
        u5_mult_82_CARRYB_43__36_), .S(u5_mult_82_SUMB_43__36_) );
  FA_X1 u5_mult_82_S2_43_35 ( .A(u5_mult_82_ab_43__35_), .B(
        u5_mult_82_CARRYB_42__35_), .CI(u5_mult_82_SUMB_42__36_), .CO(
        u5_mult_82_CARRYB_43__35_), .S(u5_mult_82_SUMB_43__35_) );
  FA_X1 u5_mult_82_S2_43_34 ( .A(u5_mult_82_ab_43__34_), .B(
        u5_mult_82_CARRYB_42__34_), .CI(u5_mult_82_SUMB_42__35_), .CO(
        u5_mult_82_CARRYB_43__34_), .S(u5_mult_82_SUMB_43__34_) );
  FA_X1 u5_mult_82_S2_43_33 ( .A(u5_mult_82_ab_43__33_), .B(
        u5_mult_82_CARRYB_42__33_), .CI(u5_mult_82_SUMB_42__34_), .CO(
        u5_mult_82_CARRYB_43__33_), .S(u5_mult_82_SUMB_43__33_) );
  FA_X1 u5_mult_82_S2_43_32 ( .A(u5_mult_82_ab_43__32_), .B(
        u5_mult_82_CARRYB_42__32_), .CI(u5_mult_82_SUMB_42__33_), .CO(
        u5_mult_82_CARRYB_43__32_), .S(u5_mult_82_SUMB_43__32_) );
  FA_X1 u5_mult_82_S2_43_31 ( .A(u5_mult_82_ab_43__31_), .B(
        u5_mult_82_CARRYB_42__31_), .CI(u5_mult_82_SUMB_42__32_), .CO(
        u5_mult_82_CARRYB_43__31_), .S(u5_mult_82_SUMB_43__31_) );
  FA_X1 u5_mult_82_S2_43_30 ( .A(u5_mult_82_ab_43__30_), .B(
        u5_mult_82_CARRYB_42__30_), .CI(u5_mult_82_SUMB_42__31_), .CO(
        u5_mult_82_CARRYB_43__30_), .S(u5_mult_82_SUMB_43__30_) );
  FA_X1 u5_mult_82_S2_43_29 ( .A(u5_mult_82_ab_43__29_), .B(
        u5_mult_82_CARRYB_42__29_), .CI(u5_mult_82_SUMB_42__30_), .CO(
        u5_mult_82_CARRYB_43__29_), .S(u5_mult_82_SUMB_43__29_) );
  FA_X1 u5_mult_82_S2_43_28 ( .A(u5_mult_82_ab_43__28_), .B(
        u5_mult_82_CARRYB_42__28_), .CI(u5_mult_82_SUMB_42__29_), .CO(
        u5_mult_82_CARRYB_43__28_), .S(u5_mult_82_SUMB_43__28_) );
  FA_X1 u5_mult_82_S2_43_27 ( .A(u5_mult_82_ab_43__27_), .B(
        u5_mult_82_CARRYB_42__27_), .CI(u5_mult_82_SUMB_42__28_), .CO(
        u5_mult_82_CARRYB_43__27_), .S(u5_mult_82_SUMB_43__27_) );
  FA_X1 u5_mult_82_S2_43_26 ( .A(u5_mult_82_ab_43__26_), .B(
        u5_mult_82_CARRYB_42__26_), .CI(u5_mult_82_SUMB_42__27_), .CO(
        u5_mult_82_CARRYB_43__26_), .S(u5_mult_82_SUMB_43__26_) );
  FA_X1 u5_mult_82_S2_43_25 ( .A(u5_mult_82_ab_43__25_), .B(
        u5_mult_82_CARRYB_42__25_), .CI(u5_mult_82_SUMB_42__26_), .CO(
        u5_mult_82_CARRYB_43__25_), .S(u5_mult_82_SUMB_43__25_) );
  FA_X1 u5_mult_82_S2_43_24 ( .A(u5_mult_82_ab_43__24_), .B(
        u5_mult_82_CARRYB_42__24_), .CI(u5_mult_82_SUMB_42__25_), .CO(
        u5_mult_82_CARRYB_43__24_), .S(u5_mult_82_SUMB_43__24_) );
  FA_X1 u5_mult_82_S2_43_23 ( .A(u5_mult_82_ab_43__23_), .B(
        u5_mult_82_CARRYB_42__23_), .CI(u5_mult_82_SUMB_42__24_), .CO(
        u5_mult_82_CARRYB_43__23_), .S(u5_mult_82_SUMB_43__23_) );
  FA_X1 u5_mult_82_S2_43_22 ( .A(u5_mult_82_ab_43__22_), .B(
        u5_mult_82_CARRYB_42__22_), .CI(u5_mult_82_SUMB_42__23_), .CO(
        u5_mult_82_CARRYB_43__22_), .S(u5_mult_82_SUMB_43__22_) );
  FA_X1 u5_mult_82_S2_43_21 ( .A(u5_mult_82_ab_43__21_), .B(
        u5_mult_82_CARRYB_42__21_), .CI(u5_mult_82_SUMB_42__22_), .CO(
        u5_mult_82_CARRYB_43__21_), .S(u5_mult_82_SUMB_43__21_) );
  FA_X1 u5_mult_82_S2_43_20 ( .A(u5_mult_82_ab_43__20_), .B(
        u5_mult_82_CARRYB_42__20_), .CI(u5_mult_82_SUMB_42__21_), .CO(
        u5_mult_82_CARRYB_43__20_), .S(u5_mult_82_SUMB_43__20_) );
  FA_X1 u5_mult_82_S2_43_19 ( .A(u5_mult_82_ab_43__19_), .B(
        u5_mult_82_CARRYB_42__19_), .CI(u5_mult_82_SUMB_42__20_), .CO(
        u5_mult_82_CARRYB_43__19_), .S(u5_mult_82_SUMB_43__19_) );
  FA_X1 u5_mult_82_S2_43_18 ( .A(u5_mult_82_ab_43__18_), .B(
        u5_mult_82_CARRYB_42__18_), .CI(u5_mult_82_SUMB_42__19_), .CO(
        u5_mult_82_CARRYB_43__18_), .S(u5_mult_82_SUMB_43__18_) );
  FA_X1 u5_mult_82_S2_43_17 ( .A(u5_mult_82_ab_43__17_), .B(
        u5_mult_82_CARRYB_42__17_), .CI(u5_mult_82_SUMB_42__18_), .CO(
        u5_mult_82_CARRYB_43__17_), .S(u5_mult_82_SUMB_43__17_) );
  FA_X1 u5_mult_82_S2_43_16 ( .A(u5_mult_82_ab_43__16_), .B(
        u5_mult_82_CARRYB_42__16_), .CI(u5_mult_82_SUMB_42__17_), .CO(
        u5_mult_82_CARRYB_43__16_), .S(u5_mult_82_SUMB_43__16_) );
  FA_X1 u5_mult_82_S2_43_15 ( .A(u5_mult_82_ab_43__15_), .B(
        u5_mult_82_CARRYB_42__15_), .CI(u5_mult_82_SUMB_42__16_), .CO(
        u5_mult_82_CARRYB_43__15_), .S(u5_mult_82_SUMB_43__15_) );
  FA_X1 u5_mult_82_S2_43_14 ( .A(u5_mult_82_ab_43__14_), .B(
        u5_mult_82_CARRYB_42__14_), .CI(u5_mult_82_SUMB_42__15_), .CO(
        u5_mult_82_CARRYB_43__14_), .S(u5_mult_82_SUMB_43__14_) );
  FA_X1 u5_mult_82_S2_43_13 ( .A(u5_mult_82_ab_43__13_), .B(
        u5_mult_82_CARRYB_42__13_), .CI(u5_mult_82_SUMB_42__14_), .CO(
        u5_mult_82_CARRYB_43__13_), .S(u5_mult_82_SUMB_43__13_) );
  FA_X1 u5_mult_82_S2_43_12 ( .A(u5_mult_82_ab_43__12_), .B(
        u5_mult_82_CARRYB_42__12_), .CI(u5_mult_82_SUMB_42__13_), .CO(
        u5_mult_82_CARRYB_43__12_), .S(u5_mult_82_SUMB_43__12_) );
  FA_X1 u5_mult_82_S2_43_11 ( .A(u5_mult_82_ab_43__11_), .B(
        u5_mult_82_CARRYB_42__11_), .CI(u5_mult_82_SUMB_42__12_), .CO(
        u5_mult_82_CARRYB_43__11_), .S(u5_mult_82_SUMB_43__11_) );
  FA_X1 u5_mult_82_S2_43_10 ( .A(u5_mult_82_ab_43__10_), .B(
        u5_mult_82_CARRYB_42__10_), .CI(u5_mult_82_SUMB_42__11_), .CO(
        u5_mult_82_CARRYB_43__10_), .S(u5_mult_82_SUMB_43__10_) );
  FA_X1 u5_mult_82_S2_43_9 ( .A(u5_mult_82_ab_43__9_), .B(
        u5_mult_82_CARRYB_42__9_), .CI(u5_mult_82_SUMB_42__10_), .CO(
        u5_mult_82_CARRYB_43__9_), .S(u5_mult_82_SUMB_43__9_) );
  FA_X1 u5_mult_82_S2_43_8 ( .A(u5_mult_82_ab_43__8_), .B(
        u5_mult_82_CARRYB_42__8_), .CI(u5_mult_82_SUMB_42__9_), .CO(
        u5_mult_82_CARRYB_43__8_), .S(u5_mult_82_SUMB_43__8_) );
  FA_X1 u5_mult_82_S2_43_7 ( .A(u5_mult_82_ab_43__7_), .B(
        u5_mult_82_CARRYB_42__7_), .CI(u5_mult_82_SUMB_42__8_), .CO(
        u5_mult_82_CARRYB_43__7_), .S(u5_mult_82_SUMB_43__7_) );
  FA_X1 u5_mult_82_S2_43_6 ( .A(u5_mult_82_ab_43__6_), .B(
        u5_mult_82_CARRYB_42__6_), .CI(u5_mult_82_SUMB_42__7_), .CO(
        u5_mult_82_CARRYB_43__6_), .S(u5_mult_82_SUMB_43__6_) );
  FA_X1 u5_mult_82_S2_43_5 ( .A(u5_mult_82_ab_43__5_), .B(
        u5_mult_82_CARRYB_42__5_), .CI(u5_mult_82_SUMB_42__6_), .CO(
        u5_mult_82_CARRYB_43__5_), .S(u5_mult_82_SUMB_43__5_) );
  FA_X1 u5_mult_82_S2_43_4 ( .A(u5_mult_82_ab_43__4_), .B(
        u5_mult_82_CARRYB_42__4_), .CI(u5_mult_82_SUMB_42__5_), .CO(
        u5_mult_82_CARRYB_43__4_), .S(u5_mult_82_SUMB_43__4_) );
  FA_X1 u5_mult_82_S2_43_3 ( .A(u5_mult_82_ab_43__3_), .B(
        u5_mult_82_CARRYB_42__3_), .CI(u5_mult_82_SUMB_42__4_), .CO(
        u5_mult_82_CARRYB_43__3_), .S(u5_mult_82_SUMB_43__3_) );
  FA_X1 u5_mult_82_S2_43_2 ( .A(u5_mult_82_ab_43__2_), .B(
        u5_mult_82_CARRYB_42__2_), .CI(u5_mult_82_SUMB_42__3_), .CO(
        u5_mult_82_CARRYB_43__2_), .S(u5_mult_82_SUMB_43__2_) );
  FA_X1 u5_mult_82_S2_43_1 ( .A(u5_mult_82_ab_43__1_), .B(
        u5_mult_82_CARRYB_42__1_), .CI(u5_mult_82_SUMB_42__2_), .CO(
        u5_mult_82_CARRYB_43__1_), .S(u5_mult_82_SUMB_43__1_) );
  FA_X1 u5_mult_82_S1_43_0 ( .A(u5_mult_82_ab_43__0_), .B(
        u5_mult_82_CARRYB_42__0_), .CI(u5_mult_82_SUMB_42__1_), .CO(
        u5_mult_82_CARRYB_43__0_), .S(u5_N43) );
  FA_X1 u5_mult_82_S3_44_51 ( .A(u5_mult_82_ab_44__51_), .B(
        u5_mult_82_CARRYB_43__51_), .CI(u5_mult_82_ab_43__52_), .CO(
        u5_mult_82_CARRYB_44__51_), .S(u5_mult_82_SUMB_44__51_) );
  FA_X1 u5_mult_82_S2_44_50 ( .A(u5_mult_82_ab_44__50_), .B(
        u5_mult_82_CARRYB_43__50_), .CI(u5_mult_82_SUMB_43__51_), .CO(
        u5_mult_82_CARRYB_44__50_), .S(u5_mult_82_SUMB_44__50_) );
  FA_X1 u5_mult_82_S2_44_49 ( .A(u5_mult_82_ab_44__49_), .B(
        u5_mult_82_CARRYB_43__49_), .CI(u5_mult_82_SUMB_43__50_), .CO(
        u5_mult_82_CARRYB_44__49_), .S(u5_mult_82_SUMB_44__49_) );
  FA_X1 u5_mult_82_S2_44_48 ( .A(u5_mult_82_ab_44__48_), .B(
        u5_mult_82_CARRYB_43__48_), .CI(u5_mult_82_SUMB_43__49_), .CO(
        u5_mult_82_CARRYB_44__48_), .S(u5_mult_82_SUMB_44__48_) );
  FA_X1 u5_mult_82_S2_44_47 ( .A(u5_mult_82_ab_44__47_), .B(
        u5_mult_82_CARRYB_43__47_), .CI(u5_mult_82_SUMB_43__48_), .CO(
        u5_mult_82_CARRYB_44__47_), .S(u5_mult_82_SUMB_44__47_) );
  FA_X1 u5_mult_82_S2_44_46 ( .A(u5_mult_82_ab_44__46_), .B(
        u5_mult_82_CARRYB_43__46_), .CI(u5_mult_82_SUMB_43__47_), .CO(
        u5_mult_82_CARRYB_44__46_), .S(u5_mult_82_SUMB_44__46_) );
  FA_X1 u5_mult_82_S2_44_45 ( .A(u5_mult_82_ab_44__45_), .B(
        u5_mult_82_CARRYB_43__45_), .CI(u5_mult_82_SUMB_43__46_), .CO(
        u5_mult_82_CARRYB_44__45_), .S(u5_mult_82_SUMB_44__45_) );
  FA_X1 u5_mult_82_S2_44_44 ( .A(u5_mult_82_ab_44__44_), .B(
        u5_mult_82_CARRYB_43__44_), .CI(u5_mult_82_SUMB_43__45_), .CO(
        u5_mult_82_CARRYB_44__44_), .S(u5_mult_82_SUMB_44__44_) );
  FA_X1 u5_mult_82_S2_44_43 ( .A(u5_mult_82_ab_44__43_), .B(
        u5_mult_82_CARRYB_43__43_), .CI(u5_mult_82_SUMB_43__44_), .CO(
        u5_mult_82_CARRYB_44__43_), .S(u5_mult_82_SUMB_44__43_) );
  FA_X1 u5_mult_82_S2_44_42 ( .A(u5_mult_82_ab_44__42_), .B(
        u5_mult_82_CARRYB_43__42_), .CI(u5_mult_82_SUMB_43__43_), .CO(
        u5_mult_82_CARRYB_44__42_), .S(u5_mult_82_SUMB_44__42_) );
  FA_X1 u5_mult_82_S2_44_41 ( .A(u5_mult_82_ab_44__41_), .B(
        u5_mult_82_CARRYB_43__41_), .CI(u5_mult_82_SUMB_43__42_), .CO(
        u5_mult_82_CARRYB_44__41_), .S(u5_mult_82_SUMB_44__41_) );
  FA_X1 u5_mult_82_S2_44_40 ( .A(u5_mult_82_ab_44__40_), .B(
        u5_mult_82_CARRYB_43__40_), .CI(u5_mult_82_SUMB_43__41_), .CO(
        u5_mult_82_CARRYB_44__40_), .S(u5_mult_82_SUMB_44__40_) );
  FA_X1 u5_mult_82_S2_44_39 ( .A(u5_mult_82_ab_44__39_), .B(
        u5_mult_82_CARRYB_43__39_), .CI(u5_mult_82_SUMB_43__40_), .CO(
        u5_mult_82_CARRYB_44__39_), .S(u5_mult_82_SUMB_44__39_) );
  FA_X1 u5_mult_82_S2_44_38 ( .A(u5_mult_82_ab_44__38_), .B(
        u5_mult_82_CARRYB_43__38_), .CI(u5_mult_82_SUMB_43__39_), .CO(
        u5_mult_82_CARRYB_44__38_), .S(u5_mult_82_SUMB_44__38_) );
  FA_X1 u5_mult_82_S2_44_37 ( .A(u5_mult_82_ab_44__37_), .B(
        u5_mult_82_CARRYB_43__37_), .CI(u5_mult_82_SUMB_43__38_), .CO(
        u5_mult_82_CARRYB_44__37_), .S(u5_mult_82_SUMB_44__37_) );
  FA_X1 u5_mult_82_S2_44_36 ( .A(u5_mult_82_ab_44__36_), .B(
        u5_mult_82_CARRYB_43__36_), .CI(u5_mult_82_SUMB_43__37_), .CO(
        u5_mult_82_CARRYB_44__36_), .S(u5_mult_82_SUMB_44__36_) );
  FA_X1 u5_mult_82_S2_44_35 ( .A(u5_mult_82_ab_44__35_), .B(
        u5_mult_82_CARRYB_43__35_), .CI(u5_mult_82_SUMB_43__36_), .CO(
        u5_mult_82_CARRYB_44__35_), .S(u5_mult_82_SUMB_44__35_) );
  FA_X1 u5_mult_82_S2_44_34 ( .A(u5_mult_82_ab_44__34_), .B(
        u5_mult_82_CARRYB_43__34_), .CI(u5_mult_82_SUMB_43__35_), .CO(
        u5_mult_82_CARRYB_44__34_), .S(u5_mult_82_SUMB_44__34_) );
  FA_X1 u5_mult_82_S2_44_33 ( .A(u5_mult_82_ab_44__33_), .B(
        u5_mult_82_CARRYB_43__33_), .CI(u5_mult_82_SUMB_43__34_), .CO(
        u5_mult_82_CARRYB_44__33_), .S(u5_mult_82_SUMB_44__33_) );
  FA_X1 u5_mult_82_S2_44_32 ( .A(u5_mult_82_ab_44__32_), .B(
        u5_mult_82_CARRYB_43__32_), .CI(u5_mult_82_SUMB_43__33_), .CO(
        u5_mult_82_CARRYB_44__32_), .S(u5_mult_82_SUMB_44__32_) );
  FA_X1 u5_mult_82_S2_44_31 ( .A(u5_mult_82_ab_44__31_), .B(
        u5_mult_82_CARRYB_43__31_), .CI(u5_mult_82_SUMB_43__32_), .CO(
        u5_mult_82_CARRYB_44__31_), .S(u5_mult_82_SUMB_44__31_) );
  FA_X1 u5_mult_82_S2_44_30 ( .A(u5_mult_82_ab_44__30_), .B(
        u5_mult_82_CARRYB_43__30_), .CI(u5_mult_82_SUMB_43__31_), .CO(
        u5_mult_82_CARRYB_44__30_), .S(u5_mult_82_SUMB_44__30_) );
  FA_X1 u5_mult_82_S2_44_29 ( .A(u5_mult_82_ab_44__29_), .B(
        u5_mult_82_CARRYB_43__29_), .CI(u5_mult_82_SUMB_43__30_), .CO(
        u5_mult_82_CARRYB_44__29_), .S(u5_mult_82_SUMB_44__29_) );
  FA_X1 u5_mult_82_S2_44_28 ( .A(u5_mult_82_ab_44__28_), .B(
        u5_mult_82_CARRYB_43__28_), .CI(u5_mult_82_SUMB_43__29_), .CO(
        u5_mult_82_CARRYB_44__28_), .S(u5_mult_82_SUMB_44__28_) );
  FA_X1 u5_mult_82_S2_44_27 ( .A(u5_mult_82_ab_44__27_), .B(
        u5_mult_82_CARRYB_43__27_), .CI(u5_mult_82_SUMB_43__28_), .CO(
        u5_mult_82_CARRYB_44__27_), .S(u5_mult_82_SUMB_44__27_) );
  FA_X1 u5_mult_82_S2_44_26 ( .A(u5_mult_82_ab_44__26_), .B(
        u5_mult_82_CARRYB_43__26_), .CI(u5_mult_82_SUMB_43__27_), .CO(
        u5_mult_82_CARRYB_44__26_), .S(u5_mult_82_SUMB_44__26_) );
  FA_X1 u5_mult_82_S2_44_25 ( .A(u5_mult_82_ab_44__25_), .B(
        u5_mult_82_CARRYB_43__25_), .CI(u5_mult_82_SUMB_43__26_), .CO(
        u5_mult_82_CARRYB_44__25_), .S(u5_mult_82_SUMB_44__25_) );
  FA_X1 u5_mult_82_S2_44_24 ( .A(u5_mult_82_ab_44__24_), .B(
        u5_mult_82_CARRYB_43__24_), .CI(u5_mult_82_SUMB_43__25_), .CO(
        u5_mult_82_CARRYB_44__24_), .S(u5_mult_82_SUMB_44__24_) );
  FA_X1 u5_mult_82_S2_44_23 ( .A(u5_mult_82_ab_44__23_), .B(
        u5_mult_82_CARRYB_43__23_), .CI(u5_mult_82_SUMB_43__24_), .CO(
        u5_mult_82_CARRYB_44__23_), .S(u5_mult_82_SUMB_44__23_) );
  FA_X1 u5_mult_82_S2_44_22 ( .A(u5_mult_82_ab_44__22_), .B(
        u5_mult_82_CARRYB_43__22_), .CI(u5_mult_82_SUMB_43__23_), .CO(
        u5_mult_82_CARRYB_44__22_), .S(u5_mult_82_SUMB_44__22_) );
  FA_X1 u5_mult_82_S2_44_21 ( .A(u5_mult_82_ab_44__21_), .B(
        u5_mult_82_CARRYB_43__21_), .CI(u5_mult_82_SUMB_43__22_), .CO(
        u5_mult_82_CARRYB_44__21_), .S(u5_mult_82_SUMB_44__21_) );
  FA_X1 u5_mult_82_S2_44_20 ( .A(u5_mult_82_ab_44__20_), .B(
        u5_mult_82_CARRYB_43__20_), .CI(u5_mult_82_SUMB_43__21_), .CO(
        u5_mult_82_CARRYB_44__20_), .S(u5_mult_82_SUMB_44__20_) );
  FA_X1 u5_mult_82_S2_44_19 ( .A(u5_mult_82_ab_44__19_), .B(
        u5_mult_82_CARRYB_43__19_), .CI(u5_mult_82_SUMB_43__20_), .CO(
        u5_mult_82_CARRYB_44__19_), .S(u5_mult_82_SUMB_44__19_) );
  FA_X1 u5_mult_82_S2_44_18 ( .A(u5_mult_82_ab_44__18_), .B(
        u5_mult_82_CARRYB_43__18_), .CI(u5_mult_82_SUMB_43__19_), .CO(
        u5_mult_82_CARRYB_44__18_), .S(u5_mult_82_SUMB_44__18_) );
  FA_X1 u5_mult_82_S2_44_17 ( .A(u5_mult_82_ab_44__17_), .B(
        u5_mult_82_CARRYB_43__17_), .CI(u5_mult_82_SUMB_43__18_), .CO(
        u5_mult_82_CARRYB_44__17_), .S(u5_mult_82_SUMB_44__17_) );
  FA_X1 u5_mult_82_S2_44_16 ( .A(u5_mult_82_ab_44__16_), .B(
        u5_mult_82_CARRYB_43__16_), .CI(u5_mult_82_SUMB_43__17_), .CO(
        u5_mult_82_CARRYB_44__16_), .S(u5_mult_82_SUMB_44__16_) );
  FA_X1 u5_mult_82_S2_44_15 ( .A(u5_mult_82_ab_44__15_), .B(
        u5_mult_82_CARRYB_43__15_), .CI(u5_mult_82_SUMB_43__16_), .CO(
        u5_mult_82_CARRYB_44__15_), .S(u5_mult_82_SUMB_44__15_) );
  FA_X1 u5_mult_82_S2_44_14 ( .A(u5_mult_82_ab_44__14_), .B(
        u5_mult_82_CARRYB_43__14_), .CI(u5_mult_82_SUMB_43__15_), .CO(
        u5_mult_82_CARRYB_44__14_), .S(u5_mult_82_SUMB_44__14_) );
  FA_X1 u5_mult_82_S2_44_13 ( .A(u5_mult_82_ab_44__13_), .B(
        u5_mult_82_CARRYB_43__13_), .CI(u5_mult_82_SUMB_43__14_), .CO(
        u5_mult_82_CARRYB_44__13_), .S(u5_mult_82_SUMB_44__13_) );
  FA_X1 u5_mult_82_S2_44_12 ( .A(u5_mult_82_ab_44__12_), .B(
        u5_mult_82_CARRYB_43__12_), .CI(u5_mult_82_SUMB_43__13_), .CO(
        u5_mult_82_CARRYB_44__12_), .S(u5_mult_82_SUMB_44__12_) );
  FA_X1 u5_mult_82_S2_44_11 ( .A(u5_mult_82_ab_44__11_), .B(
        u5_mult_82_CARRYB_43__11_), .CI(u5_mult_82_SUMB_43__12_), .CO(
        u5_mult_82_CARRYB_44__11_), .S(u5_mult_82_SUMB_44__11_) );
  FA_X1 u5_mult_82_S2_44_10 ( .A(u5_mult_82_ab_44__10_), .B(
        u5_mult_82_CARRYB_43__10_), .CI(u5_mult_82_SUMB_43__11_), .CO(
        u5_mult_82_CARRYB_44__10_), .S(u5_mult_82_SUMB_44__10_) );
  FA_X1 u5_mult_82_S2_44_9 ( .A(u5_mult_82_ab_44__9_), .B(
        u5_mult_82_CARRYB_43__9_), .CI(u5_mult_82_SUMB_43__10_), .CO(
        u5_mult_82_CARRYB_44__9_), .S(u5_mult_82_SUMB_44__9_) );
  FA_X1 u5_mult_82_S2_44_8 ( .A(u5_mult_82_ab_44__8_), .B(
        u5_mult_82_CARRYB_43__8_), .CI(u5_mult_82_SUMB_43__9_), .CO(
        u5_mult_82_CARRYB_44__8_), .S(u5_mult_82_SUMB_44__8_) );
  FA_X1 u5_mult_82_S2_44_7 ( .A(u5_mult_82_ab_44__7_), .B(
        u5_mult_82_CARRYB_43__7_), .CI(u5_mult_82_SUMB_43__8_), .CO(
        u5_mult_82_CARRYB_44__7_), .S(u5_mult_82_SUMB_44__7_) );
  FA_X1 u5_mult_82_S2_44_6 ( .A(u5_mult_82_ab_44__6_), .B(
        u5_mult_82_CARRYB_43__6_), .CI(u5_mult_82_SUMB_43__7_), .CO(
        u5_mult_82_CARRYB_44__6_), .S(u5_mult_82_SUMB_44__6_) );
  FA_X1 u5_mult_82_S2_44_5 ( .A(u5_mult_82_ab_44__5_), .B(
        u5_mult_82_CARRYB_43__5_), .CI(u5_mult_82_SUMB_43__6_), .CO(
        u5_mult_82_CARRYB_44__5_), .S(u5_mult_82_SUMB_44__5_) );
  FA_X1 u5_mult_82_S2_44_4 ( .A(u5_mult_82_ab_44__4_), .B(
        u5_mult_82_CARRYB_43__4_), .CI(u5_mult_82_SUMB_43__5_), .CO(
        u5_mult_82_CARRYB_44__4_), .S(u5_mult_82_SUMB_44__4_) );
  FA_X1 u5_mult_82_S2_44_3 ( .A(u5_mult_82_ab_44__3_), .B(
        u5_mult_82_CARRYB_43__3_), .CI(u5_mult_82_SUMB_43__4_), .CO(
        u5_mult_82_CARRYB_44__3_), .S(u5_mult_82_SUMB_44__3_) );
  FA_X1 u5_mult_82_S2_44_2 ( .A(u5_mult_82_ab_44__2_), .B(
        u5_mult_82_CARRYB_43__2_), .CI(u5_mult_82_SUMB_43__3_), .CO(
        u5_mult_82_CARRYB_44__2_), .S(u5_mult_82_SUMB_44__2_) );
  FA_X1 u5_mult_82_S2_44_1 ( .A(u5_mult_82_ab_44__1_), .B(
        u5_mult_82_CARRYB_43__1_), .CI(u5_mult_82_SUMB_43__2_), .CO(
        u5_mult_82_CARRYB_44__1_), .S(u5_mult_82_SUMB_44__1_) );
  FA_X1 u5_mult_82_S1_44_0 ( .A(u5_mult_82_ab_44__0_), .B(
        u5_mult_82_CARRYB_43__0_), .CI(u5_mult_82_SUMB_43__1_), .CO(
        u5_mult_82_CARRYB_44__0_), .S(u5_N44) );
  FA_X1 u5_mult_82_S3_45_51 ( .A(u5_mult_82_ab_45__51_), .B(
        u5_mult_82_CARRYB_44__51_), .CI(u5_mult_82_ab_44__52_), .CO(
        u5_mult_82_CARRYB_45__51_), .S(u5_mult_82_SUMB_45__51_) );
  FA_X1 u5_mult_82_S2_45_50 ( .A(u5_mult_82_ab_45__50_), .B(
        u5_mult_82_CARRYB_44__50_), .CI(u5_mult_82_SUMB_44__51_), .CO(
        u5_mult_82_CARRYB_45__50_), .S(u5_mult_82_SUMB_45__50_) );
  FA_X1 u5_mult_82_S2_45_49 ( .A(u5_mult_82_ab_45__49_), .B(
        u5_mult_82_CARRYB_44__49_), .CI(u5_mult_82_SUMB_44__50_), .CO(
        u5_mult_82_CARRYB_45__49_), .S(u5_mult_82_SUMB_45__49_) );
  FA_X1 u5_mult_82_S2_45_48 ( .A(u5_mult_82_ab_45__48_), .B(
        u5_mult_82_CARRYB_44__48_), .CI(u5_mult_82_SUMB_44__49_), .CO(
        u5_mult_82_CARRYB_45__48_), .S(u5_mult_82_SUMB_45__48_) );
  FA_X1 u5_mult_82_S2_45_47 ( .A(u5_mult_82_ab_45__47_), .B(
        u5_mult_82_CARRYB_44__47_), .CI(u5_mult_82_SUMB_44__48_), .CO(
        u5_mult_82_CARRYB_45__47_), .S(u5_mult_82_SUMB_45__47_) );
  FA_X1 u5_mult_82_S2_45_46 ( .A(u5_mult_82_ab_45__46_), .B(
        u5_mult_82_CARRYB_44__46_), .CI(u5_mult_82_SUMB_44__47_), .CO(
        u5_mult_82_CARRYB_45__46_), .S(u5_mult_82_SUMB_45__46_) );
  FA_X1 u5_mult_82_S2_45_45 ( .A(u5_mult_82_ab_45__45_), .B(
        u5_mult_82_CARRYB_44__45_), .CI(u5_mult_82_SUMB_44__46_), .CO(
        u5_mult_82_CARRYB_45__45_), .S(u5_mult_82_SUMB_45__45_) );
  FA_X1 u5_mult_82_S2_45_44 ( .A(u5_mult_82_ab_45__44_), .B(
        u5_mult_82_CARRYB_44__44_), .CI(u5_mult_82_SUMB_44__45_), .CO(
        u5_mult_82_CARRYB_45__44_), .S(u5_mult_82_SUMB_45__44_) );
  FA_X1 u5_mult_82_S2_45_43 ( .A(u5_mult_82_ab_45__43_), .B(
        u5_mult_82_CARRYB_44__43_), .CI(u5_mult_82_SUMB_44__44_), .CO(
        u5_mult_82_CARRYB_45__43_), .S(u5_mult_82_SUMB_45__43_) );
  FA_X1 u5_mult_82_S2_45_42 ( .A(u5_mult_82_ab_45__42_), .B(
        u5_mult_82_CARRYB_44__42_), .CI(u5_mult_82_SUMB_44__43_), .CO(
        u5_mult_82_CARRYB_45__42_), .S(u5_mult_82_SUMB_45__42_) );
  FA_X1 u5_mult_82_S2_45_41 ( .A(u5_mult_82_ab_45__41_), .B(
        u5_mult_82_CARRYB_44__41_), .CI(u5_mult_82_SUMB_44__42_), .CO(
        u5_mult_82_CARRYB_45__41_), .S(u5_mult_82_SUMB_45__41_) );
  FA_X1 u5_mult_82_S2_45_40 ( .A(u5_mult_82_ab_45__40_), .B(
        u5_mult_82_CARRYB_44__40_), .CI(u5_mult_82_SUMB_44__41_), .CO(
        u5_mult_82_CARRYB_45__40_), .S(u5_mult_82_SUMB_45__40_) );
  FA_X1 u5_mult_82_S2_45_39 ( .A(u5_mult_82_ab_45__39_), .B(
        u5_mult_82_CARRYB_44__39_), .CI(u5_mult_82_SUMB_44__40_), .CO(
        u5_mult_82_CARRYB_45__39_), .S(u5_mult_82_SUMB_45__39_) );
  FA_X1 u5_mult_82_S2_45_38 ( .A(u5_mult_82_ab_45__38_), .B(
        u5_mult_82_CARRYB_44__38_), .CI(u5_mult_82_SUMB_44__39_), .CO(
        u5_mult_82_CARRYB_45__38_), .S(u5_mult_82_SUMB_45__38_) );
  FA_X1 u5_mult_82_S2_45_37 ( .A(u5_mult_82_ab_45__37_), .B(
        u5_mult_82_CARRYB_44__37_), .CI(u5_mult_82_SUMB_44__38_), .CO(
        u5_mult_82_CARRYB_45__37_), .S(u5_mult_82_SUMB_45__37_) );
  FA_X1 u5_mult_82_S2_45_36 ( .A(u5_mult_82_ab_45__36_), .B(
        u5_mult_82_CARRYB_44__36_), .CI(u5_mult_82_SUMB_44__37_), .CO(
        u5_mult_82_CARRYB_45__36_), .S(u5_mult_82_SUMB_45__36_) );
  FA_X1 u5_mult_82_S2_45_35 ( .A(u5_mult_82_ab_45__35_), .B(
        u5_mult_82_CARRYB_44__35_), .CI(u5_mult_82_SUMB_44__36_), .CO(
        u5_mult_82_CARRYB_45__35_), .S(u5_mult_82_SUMB_45__35_) );
  FA_X1 u5_mult_82_S2_45_34 ( .A(u5_mult_82_ab_45__34_), .B(
        u5_mult_82_CARRYB_44__34_), .CI(u5_mult_82_SUMB_44__35_), .CO(
        u5_mult_82_CARRYB_45__34_), .S(u5_mult_82_SUMB_45__34_) );
  FA_X1 u5_mult_82_S2_45_33 ( .A(u5_mult_82_ab_45__33_), .B(
        u5_mult_82_CARRYB_44__33_), .CI(u5_mult_82_SUMB_44__34_), .CO(
        u5_mult_82_CARRYB_45__33_), .S(u5_mult_82_SUMB_45__33_) );
  FA_X1 u5_mult_82_S2_45_32 ( .A(u5_mult_82_ab_45__32_), .B(
        u5_mult_82_CARRYB_44__32_), .CI(u5_mult_82_SUMB_44__33_), .CO(
        u5_mult_82_CARRYB_45__32_), .S(u5_mult_82_SUMB_45__32_) );
  FA_X1 u5_mult_82_S2_45_31 ( .A(u5_mult_82_ab_45__31_), .B(
        u5_mult_82_CARRYB_44__31_), .CI(u5_mult_82_SUMB_44__32_), .CO(
        u5_mult_82_CARRYB_45__31_), .S(u5_mult_82_SUMB_45__31_) );
  FA_X1 u5_mult_82_S2_45_30 ( .A(u5_mult_82_ab_45__30_), .B(
        u5_mult_82_CARRYB_44__30_), .CI(u5_mult_82_SUMB_44__31_), .CO(
        u5_mult_82_CARRYB_45__30_), .S(u5_mult_82_SUMB_45__30_) );
  FA_X1 u5_mult_82_S2_45_29 ( .A(u5_mult_82_ab_45__29_), .B(
        u5_mult_82_CARRYB_44__29_), .CI(u5_mult_82_SUMB_44__30_), .CO(
        u5_mult_82_CARRYB_45__29_), .S(u5_mult_82_SUMB_45__29_) );
  FA_X1 u5_mult_82_S2_45_28 ( .A(u5_mult_82_ab_45__28_), .B(
        u5_mult_82_CARRYB_44__28_), .CI(u5_mult_82_SUMB_44__29_), .CO(
        u5_mult_82_CARRYB_45__28_), .S(u5_mult_82_SUMB_45__28_) );
  FA_X1 u5_mult_82_S2_45_27 ( .A(u5_mult_82_ab_45__27_), .B(
        u5_mult_82_CARRYB_44__27_), .CI(u5_mult_82_SUMB_44__28_), .CO(
        u5_mult_82_CARRYB_45__27_), .S(u5_mult_82_SUMB_45__27_) );
  FA_X1 u5_mult_82_S2_45_26 ( .A(u5_mult_82_ab_45__26_), .B(
        u5_mult_82_CARRYB_44__26_), .CI(u5_mult_82_SUMB_44__27_), .CO(
        u5_mult_82_CARRYB_45__26_), .S(u5_mult_82_SUMB_45__26_) );
  FA_X1 u5_mult_82_S2_45_25 ( .A(u5_mult_82_ab_45__25_), .B(
        u5_mult_82_CARRYB_44__25_), .CI(u5_mult_82_SUMB_44__26_), .CO(
        u5_mult_82_CARRYB_45__25_), .S(u5_mult_82_SUMB_45__25_) );
  FA_X1 u5_mult_82_S2_45_24 ( .A(u5_mult_82_ab_45__24_), .B(
        u5_mult_82_CARRYB_44__24_), .CI(u5_mult_82_SUMB_44__25_), .CO(
        u5_mult_82_CARRYB_45__24_), .S(u5_mult_82_SUMB_45__24_) );
  FA_X1 u5_mult_82_S2_45_23 ( .A(u5_mult_82_ab_45__23_), .B(
        u5_mult_82_CARRYB_44__23_), .CI(u5_mult_82_SUMB_44__24_), .CO(
        u5_mult_82_CARRYB_45__23_), .S(u5_mult_82_SUMB_45__23_) );
  FA_X1 u5_mult_82_S2_45_22 ( .A(u5_mult_82_ab_45__22_), .B(
        u5_mult_82_CARRYB_44__22_), .CI(u5_mult_82_SUMB_44__23_), .CO(
        u5_mult_82_CARRYB_45__22_), .S(u5_mult_82_SUMB_45__22_) );
  FA_X1 u5_mult_82_S2_45_21 ( .A(u5_mult_82_ab_45__21_), .B(
        u5_mult_82_CARRYB_44__21_), .CI(u5_mult_82_SUMB_44__22_), .CO(
        u5_mult_82_CARRYB_45__21_), .S(u5_mult_82_SUMB_45__21_) );
  FA_X1 u5_mult_82_S2_45_20 ( .A(u5_mult_82_ab_45__20_), .B(
        u5_mult_82_CARRYB_44__20_), .CI(u5_mult_82_SUMB_44__21_), .CO(
        u5_mult_82_CARRYB_45__20_), .S(u5_mult_82_SUMB_45__20_) );
  FA_X1 u5_mult_82_S2_45_19 ( .A(u5_mult_82_ab_45__19_), .B(
        u5_mult_82_CARRYB_44__19_), .CI(u5_mult_82_SUMB_44__20_), .CO(
        u5_mult_82_CARRYB_45__19_), .S(u5_mult_82_SUMB_45__19_) );
  FA_X1 u5_mult_82_S2_45_18 ( .A(u5_mult_82_ab_45__18_), .B(
        u5_mult_82_CARRYB_44__18_), .CI(u5_mult_82_SUMB_44__19_), .CO(
        u5_mult_82_CARRYB_45__18_), .S(u5_mult_82_SUMB_45__18_) );
  FA_X1 u5_mult_82_S2_45_17 ( .A(u5_mult_82_ab_45__17_), .B(
        u5_mult_82_CARRYB_44__17_), .CI(u5_mult_82_SUMB_44__18_), .CO(
        u5_mult_82_CARRYB_45__17_), .S(u5_mult_82_SUMB_45__17_) );
  FA_X1 u5_mult_82_S2_45_16 ( .A(u5_mult_82_ab_45__16_), .B(
        u5_mult_82_CARRYB_44__16_), .CI(u5_mult_82_SUMB_44__17_), .CO(
        u5_mult_82_CARRYB_45__16_), .S(u5_mult_82_SUMB_45__16_) );
  FA_X1 u5_mult_82_S2_45_15 ( .A(u5_mult_82_ab_45__15_), .B(
        u5_mult_82_CARRYB_44__15_), .CI(u5_mult_82_SUMB_44__16_), .CO(
        u5_mult_82_CARRYB_45__15_), .S(u5_mult_82_SUMB_45__15_) );
  FA_X1 u5_mult_82_S2_45_14 ( .A(u5_mult_82_ab_45__14_), .B(
        u5_mult_82_CARRYB_44__14_), .CI(u5_mult_82_SUMB_44__15_), .CO(
        u5_mult_82_CARRYB_45__14_), .S(u5_mult_82_SUMB_45__14_) );
  FA_X1 u5_mult_82_S2_45_13 ( .A(u5_mult_82_ab_45__13_), .B(
        u5_mult_82_CARRYB_44__13_), .CI(u5_mult_82_SUMB_44__14_), .CO(
        u5_mult_82_CARRYB_45__13_), .S(u5_mult_82_SUMB_45__13_) );
  FA_X1 u5_mult_82_S2_45_12 ( .A(u5_mult_82_ab_45__12_), .B(
        u5_mult_82_CARRYB_44__12_), .CI(u5_mult_82_SUMB_44__13_), .CO(
        u5_mult_82_CARRYB_45__12_), .S(u5_mult_82_SUMB_45__12_) );
  FA_X1 u5_mult_82_S2_45_11 ( .A(u5_mult_82_ab_45__11_), .B(
        u5_mult_82_CARRYB_44__11_), .CI(u5_mult_82_SUMB_44__12_), .CO(
        u5_mult_82_CARRYB_45__11_), .S(u5_mult_82_SUMB_45__11_) );
  FA_X1 u5_mult_82_S2_45_10 ( .A(u5_mult_82_ab_45__10_), .B(
        u5_mult_82_CARRYB_44__10_), .CI(u5_mult_82_SUMB_44__11_), .CO(
        u5_mult_82_CARRYB_45__10_), .S(u5_mult_82_SUMB_45__10_) );
  FA_X1 u5_mult_82_S2_45_9 ( .A(u5_mult_82_ab_45__9_), .B(
        u5_mult_82_CARRYB_44__9_), .CI(u5_mult_82_SUMB_44__10_), .CO(
        u5_mult_82_CARRYB_45__9_), .S(u5_mult_82_SUMB_45__9_) );
  FA_X1 u5_mult_82_S2_45_8 ( .A(u5_mult_82_ab_45__8_), .B(
        u5_mult_82_CARRYB_44__8_), .CI(u5_mult_82_SUMB_44__9_), .CO(
        u5_mult_82_CARRYB_45__8_), .S(u5_mult_82_SUMB_45__8_) );
  FA_X1 u5_mult_82_S2_45_7 ( .A(u5_mult_82_ab_45__7_), .B(
        u5_mult_82_CARRYB_44__7_), .CI(u5_mult_82_SUMB_44__8_), .CO(
        u5_mult_82_CARRYB_45__7_), .S(u5_mult_82_SUMB_45__7_) );
  FA_X1 u5_mult_82_S2_45_6 ( .A(u5_mult_82_ab_45__6_), .B(
        u5_mult_82_CARRYB_44__6_), .CI(u5_mult_82_SUMB_44__7_), .CO(
        u5_mult_82_CARRYB_45__6_), .S(u5_mult_82_SUMB_45__6_) );
  FA_X1 u5_mult_82_S2_45_5 ( .A(u5_mult_82_ab_45__5_), .B(
        u5_mult_82_CARRYB_44__5_), .CI(u5_mult_82_SUMB_44__6_), .CO(
        u5_mult_82_CARRYB_45__5_), .S(u5_mult_82_SUMB_45__5_) );
  FA_X1 u5_mult_82_S2_45_4 ( .A(u5_mult_82_ab_45__4_), .B(
        u5_mult_82_CARRYB_44__4_), .CI(u5_mult_82_SUMB_44__5_), .CO(
        u5_mult_82_CARRYB_45__4_), .S(u5_mult_82_SUMB_45__4_) );
  FA_X1 u5_mult_82_S2_45_3 ( .A(u5_mult_82_ab_45__3_), .B(
        u5_mult_82_CARRYB_44__3_), .CI(u5_mult_82_SUMB_44__4_), .CO(
        u5_mult_82_CARRYB_45__3_), .S(u5_mult_82_SUMB_45__3_) );
  FA_X1 u5_mult_82_S2_45_2 ( .A(u5_mult_82_ab_45__2_), .B(
        u5_mult_82_CARRYB_44__2_), .CI(u5_mult_82_SUMB_44__3_), .CO(
        u5_mult_82_CARRYB_45__2_), .S(u5_mult_82_SUMB_45__2_) );
  FA_X1 u5_mult_82_S2_45_1 ( .A(u5_mult_82_ab_45__1_), .B(
        u5_mult_82_CARRYB_44__1_), .CI(u5_mult_82_SUMB_44__2_), .CO(
        u5_mult_82_CARRYB_45__1_), .S(u5_mult_82_SUMB_45__1_) );
  FA_X1 u5_mult_82_S1_45_0 ( .A(u5_mult_82_ab_45__0_), .B(
        u5_mult_82_CARRYB_44__0_), .CI(u5_mult_82_SUMB_44__1_), .CO(
        u5_mult_82_CARRYB_45__0_), .S(u5_N45) );
  FA_X1 u5_mult_82_S3_46_51 ( .A(u5_mult_82_ab_46__51_), .B(
        u5_mult_82_CARRYB_45__51_), .CI(u5_mult_82_ab_45__52_), .CO(
        u5_mult_82_CARRYB_46__51_), .S(u5_mult_82_SUMB_46__51_) );
  FA_X1 u5_mult_82_S2_46_50 ( .A(u5_mult_82_ab_46__50_), .B(
        u5_mult_82_CARRYB_45__50_), .CI(u5_mult_82_SUMB_45__51_), .CO(
        u5_mult_82_CARRYB_46__50_), .S(u5_mult_82_SUMB_46__50_) );
  FA_X1 u5_mult_82_S2_46_49 ( .A(u5_mult_82_ab_46__49_), .B(
        u5_mult_82_CARRYB_45__49_), .CI(u5_mult_82_SUMB_45__50_), .CO(
        u5_mult_82_CARRYB_46__49_), .S(u5_mult_82_SUMB_46__49_) );
  FA_X1 u5_mult_82_S2_46_48 ( .A(u5_mult_82_ab_46__48_), .B(
        u5_mult_82_CARRYB_45__48_), .CI(u5_mult_82_SUMB_45__49_), .CO(
        u5_mult_82_CARRYB_46__48_), .S(u5_mult_82_SUMB_46__48_) );
  FA_X1 u5_mult_82_S2_46_47 ( .A(u5_mult_82_ab_46__47_), .B(
        u5_mult_82_CARRYB_45__47_), .CI(u5_mult_82_SUMB_45__48_), .CO(
        u5_mult_82_CARRYB_46__47_), .S(u5_mult_82_SUMB_46__47_) );
  FA_X1 u5_mult_82_S2_46_46 ( .A(u5_mult_82_ab_46__46_), .B(
        u5_mult_82_CARRYB_45__46_), .CI(u5_mult_82_SUMB_45__47_), .CO(
        u5_mult_82_CARRYB_46__46_), .S(u5_mult_82_SUMB_46__46_) );
  FA_X1 u5_mult_82_S2_46_45 ( .A(u5_mult_82_ab_46__45_), .B(
        u5_mult_82_CARRYB_45__45_), .CI(u5_mult_82_SUMB_45__46_), .CO(
        u5_mult_82_CARRYB_46__45_), .S(u5_mult_82_SUMB_46__45_) );
  FA_X1 u5_mult_82_S2_46_44 ( .A(u5_mult_82_ab_46__44_), .B(
        u5_mult_82_CARRYB_45__44_), .CI(u5_mult_82_SUMB_45__45_), .CO(
        u5_mult_82_CARRYB_46__44_), .S(u5_mult_82_SUMB_46__44_) );
  FA_X1 u5_mult_82_S2_46_43 ( .A(u5_mult_82_ab_46__43_), .B(
        u5_mult_82_CARRYB_45__43_), .CI(u5_mult_82_SUMB_45__44_), .CO(
        u5_mult_82_CARRYB_46__43_), .S(u5_mult_82_SUMB_46__43_) );
  FA_X1 u5_mult_82_S2_46_42 ( .A(u5_mult_82_ab_46__42_), .B(
        u5_mult_82_CARRYB_45__42_), .CI(u5_mult_82_SUMB_45__43_), .CO(
        u5_mult_82_CARRYB_46__42_), .S(u5_mult_82_SUMB_46__42_) );
  FA_X1 u5_mult_82_S2_46_41 ( .A(u5_mult_82_ab_46__41_), .B(
        u5_mult_82_CARRYB_45__41_), .CI(u5_mult_82_SUMB_45__42_), .CO(
        u5_mult_82_CARRYB_46__41_), .S(u5_mult_82_SUMB_46__41_) );
  FA_X1 u5_mult_82_S2_46_40 ( .A(u5_mult_82_ab_46__40_), .B(
        u5_mult_82_CARRYB_45__40_), .CI(u5_mult_82_SUMB_45__41_), .CO(
        u5_mult_82_CARRYB_46__40_), .S(u5_mult_82_SUMB_46__40_) );
  FA_X1 u5_mult_82_S2_46_39 ( .A(u5_mult_82_ab_46__39_), .B(
        u5_mult_82_CARRYB_45__39_), .CI(u5_mult_82_SUMB_45__40_), .CO(
        u5_mult_82_CARRYB_46__39_), .S(u5_mult_82_SUMB_46__39_) );
  FA_X1 u5_mult_82_S2_46_38 ( .A(u5_mult_82_ab_46__38_), .B(
        u5_mult_82_CARRYB_45__38_), .CI(u5_mult_82_SUMB_45__39_), .CO(
        u5_mult_82_CARRYB_46__38_), .S(u5_mult_82_SUMB_46__38_) );
  FA_X1 u5_mult_82_S2_46_37 ( .A(u5_mult_82_ab_46__37_), .B(
        u5_mult_82_CARRYB_45__37_), .CI(u5_mult_82_SUMB_45__38_), .CO(
        u5_mult_82_CARRYB_46__37_), .S(u5_mult_82_SUMB_46__37_) );
  FA_X1 u5_mult_82_S2_46_36 ( .A(u5_mult_82_ab_46__36_), .B(
        u5_mult_82_CARRYB_45__36_), .CI(u5_mult_82_SUMB_45__37_), .CO(
        u5_mult_82_CARRYB_46__36_), .S(u5_mult_82_SUMB_46__36_) );
  FA_X1 u5_mult_82_S2_46_35 ( .A(u5_mult_82_ab_46__35_), .B(
        u5_mult_82_CARRYB_45__35_), .CI(u5_mult_82_SUMB_45__36_), .CO(
        u5_mult_82_CARRYB_46__35_), .S(u5_mult_82_SUMB_46__35_) );
  FA_X1 u5_mult_82_S2_46_34 ( .A(u5_mult_82_ab_46__34_), .B(
        u5_mult_82_CARRYB_45__34_), .CI(u5_mult_82_SUMB_45__35_), .CO(
        u5_mult_82_CARRYB_46__34_), .S(u5_mult_82_SUMB_46__34_) );
  FA_X1 u5_mult_82_S2_46_33 ( .A(u5_mult_82_ab_46__33_), .B(
        u5_mult_82_CARRYB_45__33_), .CI(u5_mult_82_SUMB_45__34_), .CO(
        u5_mult_82_CARRYB_46__33_), .S(u5_mult_82_SUMB_46__33_) );
  FA_X1 u5_mult_82_S2_46_32 ( .A(u5_mult_82_ab_46__32_), .B(
        u5_mult_82_CARRYB_45__32_), .CI(u5_mult_82_SUMB_45__33_), .CO(
        u5_mult_82_CARRYB_46__32_), .S(u5_mult_82_SUMB_46__32_) );
  FA_X1 u5_mult_82_S2_46_31 ( .A(u5_mult_82_ab_46__31_), .B(
        u5_mult_82_CARRYB_45__31_), .CI(u5_mult_82_SUMB_45__32_), .CO(
        u5_mult_82_CARRYB_46__31_), .S(u5_mult_82_SUMB_46__31_) );
  FA_X1 u5_mult_82_S2_46_30 ( .A(u5_mult_82_ab_46__30_), .B(
        u5_mult_82_CARRYB_45__30_), .CI(u5_mult_82_SUMB_45__31_), .CO(
        u5_mult_82_CARRYB_46__30_), .S(u5_mult_82_SUMB_46__30_) );
  FA_X1 u5_mult_82_S2_46_29 ( .A(u5_mult_82_ab_46__29_), .B(
        u5_mult_82_CARRYB_45__29_), .CI(u5_mult_82_SUMB_45__30_), .CO(
        u5_mult_82_CARRYB_46__29_), .S(u5_mult_82_SUMB_46__29_) );
  FA_X1 u5_mult_82_S2_46_28 ( .A(u5_mult_82_ab_46__28_), .B(
        u5_mult_82_CARRYB_45__28_), .CI(u5_mult_82_SUMB_45__29_), .CO(
        u5_mult_82_CARRYB_46__28_), .S(u5_mult_82_SUMB_46__28_) );
  FA_X1 u5_mult_82_S2_46_27 ( .A(u5_mult_82_ab_46__27_), .B(
        u5_mult_82_CARRYB_45__27_), .CI(u5_mult_82_SUMB_45__28_), .CO(
        u5_mult_82_CARRYB_46__27_), .S(u5_mult_82_SUMB_46__27_) );
  FA_X1 u5_mult_82_S2_46_26 ( .A(u5_mult_82_ab_46__26_), .B(
        u5_mult_82_CARRYB_45__26_), .CI(u5_mult_82_SUMB_45__27_), .CO(
        u5_mult_82_CARRYB_46__26_), .S(u5_mult_82_SUMB_46__26_) );
  FA_X1 u5_mult_82_S2_46_25 ( .A(u5_mult_82_ab_46__25_), .B(
        u5_mult_82_CARRYB_45__25_), .CI(u5_mult_82_SUMB_45__26_), .CO(
        u5_mult_82_CARRYB_46__25_), .S(u5_mult_82_SUMB_46__25_) );
  FA_X1 u5_mult_82_S2_46_24 ( .A(u5_mult_82_ab_46__24_), .B(
        u5_mult_82_CARRYB_45__24_), .CI(u5_mult_82_SUMB_45__25_), .CO(
        u5_mult_82_CARRYB_46__24_), .S(u5_mult_82_SUMB_46__24_) );
  FA_X1 u5_mult_82_S2_46_23 ( .A(u5_mult_82_ab_46__23_), .B(
        u5_mult_82_CARRYB_45__23_), .CI(u5_mult_82_SUMB_45__24_), .CO(
        u5_mult_82_CARRYB_46__23_), .S(u5_mult_82_SUMB_46__23_) );
  FA_X1 u5_mult_82_S2_46_22 ( .A(u5_mult_82_ab_46__22_), .B(
        u5_mult_82_CARRYB_45__22_), .CI(u5_mult_82_SUMB_45__23_), .CO(
        u5_mult_82_CARRYB_46__22_), .S(u5_mult_82_SUMB_46__22_) );
  FA_X1 u5_mult_82_S2_46_21 ( .A(u5_mult_82_ab_46__21_), .B(
        u5_mult_82_CARRYB_45__21_), .CI(u5_mult_82_SUMB_45__22_), .CO(
        u5_mult_82_CARRYB_46__21_), .S(u5_mult_82_SUMB_46__21_) );
  FA_X1 u5_mult_82_S2_46_20 ( .A(u5_mult_82_ab_46__20_), .B(
        u5_mult_82_CARRYB_45__20_), .CI(u5_mult_82_SUMB_45__21_), .CO(
        u5_mult_82_CARRYB_46__20_), .S(u5_mult_82_SUMB_46__20_) );
  FA_X1 u5_mult_82_S2_46_19 ( .A(u5_mult_82_ab_46__19_), .B(
        u5_mult_82_CARRYB_45__19_), .CI(u5_mult_82_SUMB_45__20_), .CO(
        u5_mult_82_CARRYB_46__19_), .S(u5_mult_82_SUMB_46__19_) );
  FA_X1 u5_mult_82_S2_46_18 ( .A(u5_mult_82_ab_46__18_), .B(
        u5_mult_82_CARRYB_45__18_), .CI(u5_mult_82_SUMB_45__19_), .CO(
        u5_mult_82_CARRYB_46__18_), .S(u5_mult_82_SUMB_46__18_) );
  FA_X1 u5_mult_82_S2_46_17 ( .A(u5_mult_82_ab_46__17_), .B(
        u5_mult_82_CARRYB_45__17_), .CI(u5_mult_82_SUMB_45__18_), .CO(
        u5_mult_82_CARRYB_46__17_), .S(u5_mult_82_SUMB_46__17_) );
  FA_X1 u5_mult_82_S2_46_16 ( .A(u5_mult_82_ab_46__16_), .B(
        u5_mult_82_CARRYB_45__16_), .CI(u5_mult_82_SUMB_45__17_), .CO(
        u5_mult_82_CARRYB_46__16_), .S(u5_mult_82_SUMB_46__16_) );
  FA_X1 u5_mult_82_S2_46_15 ( .A(u5_mult_82_ab_46__15_), .B(
        u5_mult_82_CARRYB_45__15_), .CI(u5_mult_82_SUMB_45__16_), .CO(
        u5_mult_82_CARRYB_46__15_), .S(u5_mult_82_SUMB_46__15_) );
  FA_X1 u5_mult_82_S2_46_14 ( .A(u5_mult_82_ab_46__14_), .B(
        u5_mult_82_CARRYB_45__14_), .CI(u5_mult_82_SUMB_45__15_), .CO(
        u5_mult_82_CARRYB_46__14_), .S(u5_mult_82_SUMB_46__14_) );
  FA_X1 u5_mult_82_S2_46_13 ( .A(u5_mult_82_ab_46__13_), .B(
        u5_mult_82_CARRYB_45__13_), .CI(u5_mult_82_SUMB_45__14_), .CO(
        u5_mult_82_CARRYB_46__13_), .S(u5_mult_82_SUMB_46__13_) );
  FA_X1 u5_mult_82_S2_46_12 ( .A(u5_mult_82_ab_46__12_), .B(
        u5_mult_82_CARRYB_45__12_), .CI(u5_mult_82_SUMB_45__13_), .CO(
        u5_mult_82_CARRYB_46__12_), .S(u5_mult_82_SUMB_46__12_) );
  FA_X1 u5_mult_82_S2_46_11 ( .A(u5_mult_82_ab_46__11_), .B(
        u5_mult_82_CARRYB_45__11_), .CI(u5_mult_82_SUMB_45__12_), .CO(
        u5_mult_82_CARRYB_46__11_), .S(u5_mult_82_SUMB_46__11_) );
  FA_X1 u5_mult_82_S2_46_10 ( .A(u5_mult_82_ab_46__10_), .B(
        u5_mult_82_CARRYB_45__10_), .CI(u5_mult_82_SUMB_45__11_), .CO(
        u5_mult_82_CARRYB_46__10_), .S(u5_mult_82_SUMB_46__10_) );
  FA_X1 u5_mult_82_S2_46_9 ( .A(u5_mult_82_ab_46__9_), .B(
        u5_mult_82_CARRYB_45__9_), .CI(u5_mult_82_SUMB_45__10_), .CO(
        u5_mult_82_CARRYB_46__9_), .S(u5_mult_82_SUMB_46__9_) );
  FA_X1 u5_mult_82_S2_46_8 ( .A(u5_mult_82_ab_46__8_), .B(
        u5_mult_82_CARRYB_45__8_), .CI(u5_mult_82_SUMB_45__9_), .CO(
        u5_mult_82_CARRYB_46__8_), .S(u5_mult_82_SUMB_46__8_) );
  FA_X1 u5_mult_82_S2_46_7 ( .A(u5_mult_82_ab_46__7_), .B(
        u5_mult_82_CARRYB_45__7_), .CI(u5_mult_82_SUMB_45__8_), .CO(
        u5_mult_82_CARRYB_46__7_), .S(u5_mult_82_SUMB_46__7_) );
  FA_X1 u5_mult_82_S2_46_6 ( .A(u5_mult_82_ab_46__6_), .B(
        u5_mult_82_CARRYB_45__6_), .CI(u5_mult_82_SUMB_45__7_), .CO(
        u5_mult_82_CARRYB_46__6_), .S(u5_mult_82_SUMB_46__6_) );
  FA_X1 u5_mult_82_S2_46_5 ( .A(u5_mult_82_ab_46__5_), .B(
        u5_mult_82_CARRYB_45__5_), .CI(u5_mult_82_SUMB_45__6_), .CO(
        u5_mult_82_CARRYB_46__5_), .S(u5_mult_82_SUMB_46__5_) );
  FA_X1 u5_mult_82_S2_46_4 ( .A(u5_mult_82_ab_46__4_), .B(
        u5_mult_82_CARRYB_45__4_), .CI(u5_mult_82_SUMB_45__5_), .CO(
        u5_mult_82_CARRYB_46__4_), .S(u5_mult_82_SUMB_46__4_) );
  FA_X1 u5_mult_82_S2_46_3 ( .A(u5_mult_82_ab_46__3_), .B(
        u5_mult_82_CARRYB_45__3_), .CI(u5_mult_82_SUMB_45__4_), .CO(
        u5_mult_82_CARRYB_46__3_), .S(u5_mult_82_SUMB_46__3_) );
  FA_X1 u5_mult_82_S2_46_2 ( .A(u5_mult_82_ab_46__2_), .B(
        u5_mult_82_CARRYB_45__2_), .CI(u5_mult_82_SUMB_45__3_), .CO(
        u5_mult_82_CARRYB_46__2_), .S(u5_mult_82_SUMB_46__2_) );
  FA_X1 u5_mult_82_S2_46_1 ( .A(u5_mult_82_ab_46__1_), .B(
        u5_mult_82_CARRYB_45__1_), .CI(u5_mult_82_SUMB_45__2_), .CO(
        u5_mult_82_CARRYB_46__1_), .S(u5_mult_82_SUMB_46__1_) );
  FA_X1 u5_mult_82_S1_46_0 ( .A(u5_mult_82_ab_46__0_), .B(
        u5_mult_82_CARRYB_45__0_), .CI(u5_mult_82_SUMB_45__1_), .CO(
        u5_mult_82_CARRYB_46__0_), .S(u5_N46) );
  FA_X1 u5_mult_82_S3_47_51 ( .A(u5_mult_82_ab_47__51_), .B(
        u5_mult_82_CARRYB_46__51_), .CI(u5_mult_82_ab_46__52_), .CO(
        u5_mult_82_CARRYB_47__51_), .S(u5_mult_82_SUMB_47__51_) );
  FA_X1 u5_mult_82_S2_47_50 ( .A(u5_mult_82_ab_47__50_), .B(
        u5_mult_82_CARRYB_46__50_), .CI(u5_mult_82_SUMB_46__51_), .CO(
        u5_mult_82_CARRYB_47__50_), .S(u5_mult_82_SUMB_47__50_) );
  FA_X1 u5_mult_82_S2_47_49 ( .A(u5_mult_82_ab_47__49_), .B(
        u5_mult_82_CARRYB_46__49_), .CI(u5_mult_82_SUMB_46__50_), .CO(
        u5_mult_82_CARRYB_47__49_), .S(u5_mult_82_SUMB_47__49_) );
  FA_X1 u5_mult_82_S2_47_48 ( .A(u5_mult_82_ab_47__48_), .B(
        u5_mult_82_CARRYB_46__48_), .CI(u5_mult_82_SUMB_46__49_), .CO(
        u5_mult_82_CARRYB_47__48_), .S(u5_mult_82_SUMB_47__48_) );
  FA_X1 u5_mult_82_S2_47_47 ( .A(u5_mult_82_ab_47__47_), .B(
        u5_mult_82_CARRYB_46__47_), .CI(u5_mult_82_SUMB_46__48_), .CO(
        u5_mult_82_CARRYB_47__47_), .S(u5_mult_82_SUMB_47__47_) );
  FA_X1 u5_mult_82_S2_47_46 ( .A(u5_mult_82_ab_47__46_), .B(
        u5_mult_82_CARRYB_46__46_), .CI(u5_mult_82_SUMB_46__47_), .CO(
        u5_mult_82_CARRYB_47__46_), .S(u5_mult_82_SUMB_47__46_) );
  FA_X1 u5_mult_82_S2_47_45 ( .A(u5_mult_82_ab_47__45_), .B(
        u5_mult_82_CARRYB_46__45_), .CI(u5_mult_82_SUMB_46__46_), .CO(
        u5_mult_82_CARRYB_47__45_), .S(u5_mult_82_SUMB_47__45_) );
  FA_X1 u5_mult_82_S2_47_44 ( .A(u5_mult_82_ab_47__44_), .B(
        u5_mult_82_CARRYB_46__44_), .CI(u5_mult_82_SUMB_46__45_), .CO(
        u5_mult_82_CARRYB_47__44_), .S(u5_mult_82_SUMB_47__44_) );
  FA_X1 u5_mult_82_S2_47_43 ( .A(u5_mult_82_ab_47__43_), .B(
        u5_mult_82_CARRYB_46__43_), .CI(u5_mult_82_SUMB_46__44_), .CO(
        u5_mult_82_CARRYB_47__43_), .S(u5_mult_82_SUMB_47__43_) );
  FA_X1 u5_mult_82_S2_47_42 ( .A(u5_mult_82_ab_47__42_), .B(
        u5_mult_82_CARRYB_46__42_), .CI(u5_mult_82_SUMB_46__43_), .CO(
        u5_mult_82_CARRYB_47__42_), .S(u5_mult_82_SUMB_47__42_) );
  FA_X1 u5_mult_82_S2_47_41 ( .A(u5_mult_82_ab_47__41_), .B(
        u5_mult_82_CARRYB_46__41_), .CI(u5_mult_82_SUMB_46__42_), .CO(
        u5_mult_82_CARRYB_47__41_), .S(u5_mult_82_SUMB_47__41_) );
  FA_X1 u5_mult_82_S2_47_40 ( .A(u5_mult_82_ab_47__40_), .B(
        u5_mult_82_CARRYB_46__40_), .CI(u5_mult_82_SUMB_46__41_), .CO(
        u5_mult_82_CARRYB_47__40_), .S(u5_mult_82_SUMB_47__40_) );
  FA_X1 u5_mult_82_S2_47_39 ( .A(u5_mult_82_ab_47__39_), .B(
        u5_mult_82_CARRYB_46__39_), .CI(u5_mult_82_SUMB_46__40_), .CO(
        u5_mult_82_CARRYB_47__39_), .S(u5_mult_82_SUMB_47__39_) );
  FA_X1 u5_mult_82_S2_47_38 ( .A(u5_mult_82_ab_47__38_), .B(
        u5_mult_82_CARRYB_46__38_), .CI(u5_mult_82_SUMB_46__39_), .CO(
        u5_mult_82_CARRYB_47__38_), .S(u5_mult_82_SUMB_47__38_) );
  FA_X1 u5_mult_82_S2_47_37 ( .A(u5_mult_82_ab_47__37_), .B(
        u5_mult_82_CARRYB_46__37_), .CI(u5_mult_82_SUMB_46__38_), .CO(
        u5_mult_82_CARRYB_47__37_), .S(u5_mult_82_SUMB_47__37_) );
  FA_X1 u5_mult_82_S2_47_36 ( .A(u5_mult_82_ab_47__36_), .B(
        u5_mult_82_CARRYB_46__36_), .CI(u5_mult_82_SUMB_46__37_), .CO(
        u5_mult_82_CARRYB_47__36_), .S(u5_mult_82_SUMB_47__36_) );
  FA_X1 u5_mult_82_S2_47_35 ( .A(u5_mult_82_ab_47__35_), .B(
        u5_mult_82_CARRYB_46__35_), .CI(u5_mult_82_SUMB_46__36_), .CO(
        u5_mult_82_CARRYB_47__35_), .S(u5_mult_82_SUMB_47__35_) );
  FA_X1 u5_mult_82_S2_47_34 ( .A(u5_mult_82_ab_47__34_), .B(
        u5_mult_82_CARRYB_46__34_), .CI(u5_mult_82_SUMB_46__35_), .CO(
        u5_mult_82_CARRYB_47__34_), .S(u5_mult_82_SUMB_47__34_) );
  FA_X1 u5_mult_82_S2_47_33 ( .A(u5_mult_82_ab_47__33_), .B(
        u5_mult_82_CARRYB_46__33_), .CI(u5_mult_82_SUMB_46__34_), .CO(
        u5_mult_82_CARRYB_47__33_), .S(u5_mult_82_SUMB_47__33_) );
  FA_X1 u5_mult_82_S2_47_32 ( .A(u5_mult_82_ab_47__32_), .B(
        u5_mult_82_CARRYB_46__32_), .CI(u5_mult_82_SUMB_46__33_), .CO(
        u5_mult_82_CARRYB_47__32_), .S(u5_mult_82_SUMB_47__32_) );
  FA_X1 u5_mult_82_S2_47_31 ( .A(u5_mult_82_ab_47__31_), .B(
        u5_mult_82_CARRYB_46__31_), .CI(u5_mult_82_SUMB_46__32_), .CO(
        u5_mult_82_CARRYB_47__31_), .S(u5_mult_82_SUMB_47__31_) );
  FA_X1 u5_mult_82_S2_47_30 ( .A(u5_mult_82_ab_47__30_), .B(
        u5_mult_82_CARRYB_46__30_), .CI(u5_mult_82_SUMB_46__31_), .CO(
        u5_mult_82_CARRYB_47__30_), .S(u5_mult_82_SUMB_47__30_) );
  FA_X1 u5_mult_82_S2_47_29 ( .A(u5_mult_82_ab_47__29_), .B(
        u5_mult_82_CARRYB_46__29_), .CI(u5_mult_82_SUMB_46__30_), .CO(
        u5_mult_82_CARRYB_47__29_), .S(u5_mult_82_SUMB_47__29_) );
  FA_X1 u5_mult_82_S2_47_28 ( .A(u5_mult_82_ab_47__28_), .B(
        u5_mult_82_CARRYB_46__28_), .CI(u5_mult_82_SUMB_46__29_), .CO(
        u5_mult_82_CARRYB_47__28_), .S(u5_mult_82_SUMB_47__28_) );
  FA_X1 u5_mult_82_S2_47_27 ( .A(u5_mult_82_ab_47__27_), .B(
        u5_mult_82_CARRYB_46__27_), .CI(u5_mult_82_SUMB_46__28_), .CO(
        u5_mult_82_CARRYB_47__27_), .S(u5_mult_82_SUMB_47__27_) );
  FA_X1 u5_mult_82_S2_47_26 ( .A(u5_mult_82_ab_47__26_), .B(
        u5_mult_82_CARRYB_46__26_), .CI(u5_mult_82_SUMB_46__27_), .CO(
        u5_mult_82_CARRYB_47__26_), .S(u5_mult_82_SUMB_47__26_) );
  FA_X1 u5_mult_82_S2_47_25 ( .A(u5_mult_82_ab_47__25_), .B(
        u5_mult_82_CARRYB_46__25_), .CI(u5_mult_82_SUMB_46__26_), .CO(
        u5_mult_82_CARRYB_47__25_), .S(u5_mult_82_SUMB_47__25_) );
  FA_X1 u5_mult_82_S2_47_24 ( .A(u5_mult_82_ab_47__24_), .B(
        u5_mult_82_CARRYB_46__24_), .CI(u5_mult_82_SUMB_46__25_), .CO(
        u5_mult_82_CARRYB_47__24_), .S(u5_mult_82_SUMB_47__24_) );
  FA_X1 u5_mult_82_S2_47_23 ( .A(u5_mult_82_ab_47__23_), .B(
        u5_mult_82_CARRYB_46__23_), .CI(u5_mult_82_SUMB_46__24_), .CO(
        u5_mult_82_CARRYB_47__23_), .S(u5_mult_82_SUMB_47__23_) );
  FA_X1 u5_mult_82_S2_47_22 ( .A(u5_mult_82_ab_47__22_), .B(
        u5_mult_82_CARRYB_46__22_), .CI(u5_mult_82_SUMB_46__23_), .CO(
        u5_mult_82_CARRYB_47__22_), .S(u5_mult_82_SUMB_47__22_) );
  FA_X1 u5_mult_82_S2_47_21 ( .A(u5_mult_82_ab_47__21_), .B(
        u5_mult_82_CARRYB_46__21_), .CI(u5_mult_82_SUMB_46__22_), .CO(
        u5_mult_82_CARRYB_47__21_), .S(u5_mult_82_SUMB_47__21_) );
  FA_X1 u5_mult_82_S2_47_20 ( .A(u5_mult_82_ab_47__20_), .B(
        u5_mult_82_CARRYB_46__20_), .CI(u5_mult_82_SUMB_46__21_), .CO(
        u5_mult_82_CARRYB_47__20_), .S(u5_mult_82_SUMB_47__20_) );
  FA_X1 u5_mult_82_S2_47_19 ( .A(u5_mult_82_ab_47__19_), .B(
        u5_mult_82_CARRYB_46__19_), .CI(u5_mult_82_SUMB_46__20_), .CO(
        u5_mult_82_CARRYB_47__19_), .S(u5_mult_82_SUMB_47__19_) );
  FA_X1 u5_mult_82_S2_47_18 ( .A(u5_mult_82_ab_47__18_), .B(
        u5_mult_82_CARRYB_46__18_), .CI(u5_mult_82_SUMB_46__19_), .CO(
        u5_mult_82_CARRYB_47__18_), .S(u5_mult_82_SUMB_47__18_) );
  FA_X1 u5_mult_82_S2_47_17 ( .A(u5_mult_82_ab_47__17_), .B(
        u5_mult_82_CARRYB_46__17_), .CI(u5_mult_82_SUMB_46__18_), .CO(
        u5_mult_82_CARRYB_47__17_), .S(u5_mult_82_SUMB_47__17_) );
  FA_X1 u5_mult_82_S2_47_16 ( .A(u5_mult_82_ab_47__16_), .B(
        u5_mult_82_CARRYB_46__16_), .CI(u5_mult_82_SUMB_46__17_), .CO(
        u5_mult_82_CARRYB_47__16_), .S(u5_mult_82_SUMB_47__16_) );
  FA_X1 u5_mult_82_S2_47_15 ( .A(u5_mult_82_ab_47__15_), .B(
        u5_mult_82_CARRYB_46__15_), .CI(u5_mult_82_SUMB_46__16_), .CO(
        u5_mult_82_CARRYB_47__15_), .S(u5_mult_82_SUMB_47__15_) );
  FA_X1 u5_mult_82_S2_47_14 ( .A(u5_mult_82_ab_47__14_), .B(
        u5_mult_82_CARRYB_46__14_), .CI(u5_mult_82_SUMB_46__15_), .CO(
        u5_mult_82_CARRYB_47__14_), .S(u5_mult_82_SUMB_47__14_) );
  FA_X1 u5_mult_82_S2_47_13 ( .A(u5_mult_82_ab_47__13_), .B(
        u5_mult_82_CARRYB_46__13_), .CI(u5_mult_82_SUMB_46__14_), .CO(
        u5_mult_82_CARRYB_47__13_), .S(u5_mult_82_SUMB_47__13_) );
  FA_X1 u5_mult_82_S2_47_12 ( .A(u5_mult_82_ab_47__12_), .B(
        u5_mult_82_CARRYB_46__12_), .CI(u5_mult_82_SUMB_46__13_), .CO(
        u5_mult_82_CARRYB_47__12_), .S(u5_mult_82_SUMB_47__12_) );
  FA_X1 u5_mult_82_S2_47_11 ( .A(u5_mult_82_ab_47__11_), .B(
        u5_mult_82_CARRYB_46__11_), .CI(u5_mult_82_SUMB_46__12_), .CO(
        u5_mult_82_CARRYB_47__11_), .S(u5_mult_82_SUMB_47__11_) );
  FA_X1 u5_mult_82_S2_47_10 ( .A(u5_mult_82_ab_47__10_), .B(
        u5_mult_82_CARRYB_46__10_), .CI(u5_mult_82_SUMB_46__11_), .CO(
        u5_mult_82_CARRYB_47__10_), .S(u5_mult_82_SUMB_47__10_) );
  FA_X1 u5_mult_82_S2_47_9 ( .A(u5_mult_82_ab_47__9_), .B(
        u5_mult_82_CARRYB_46__9_), .CI(u5_mult_82_SUMB_46__10_), .CO(
        u5_mult_82_CARRYB_47__9_), .S(u5_mult_82_SUMB_47__9_) );
  FA_X1 u5_mult_82_S2_47_8 ( .A(u5_mult_82_ab_47__8_), .B(
        u5_mult_82_CARRYB_46__8_), .CI(u5_mult_82_SUMB_46__9_), .CO(
        u5_mult_82_CARRYB_47__8_), .S(u5_mult_82_SUMB_47__8_) );
  FA_X1 u5_mult_82_S2_47_7 ( .A(u5_mult_82_ab_47__7_), .B(
        u5_mult_82_CARRYB_46__7_), .CI(u5_mult_82_SUMB_46__8_), .CO(
        u5_mult_82_CARRYB_47__7_), .S(u5_mult_82_SUMB_47__7_) );
  FA_X1 u5_mult_82_S2_47_6 ( .A(u5_mult_82_ab_47__6_), .B(
        u5_mult_82_CARRYB_46__6_), .CI(u5_mult_82_SUMB_46__7_), .CO(
        u5_mult_82_CARRYB_47__6_), .S(u5_mult_82_SUMB_47__6_) );
  FA_X1 u5_mult_82_S2_47_5 ( .A(u5_mult_82_ab_47__5_), .B(
        u5_mult_82_CARRYB_46__5_), .CI(u5_mult_82_SUMB_46__6_), .CO(
        u5_mult_82_CARRYB_47__5_), .S(u5_mult_82_SUMB_47__5_) );
  FA_X1 u5_mult_82_S2_47_4 ( .A(u5_mult_82_ab_47__4_), .B(
        u5_mult_82_CARRYB_46__4_), .CI(u5_mult_82_SUMB_46__5_), .CO(
        u5_mult_82_CARRYB_47__4_), .S(u5_mult_82_SUMB_47__4_) );
  FA_X1 u5_mult_82_S2_47_3 ( .A(u5_mult_82_ab_47__3_), .B(
        u5_mult_82_CARRYB_46__3_), .CI(u5_mult_82_SUMB_46__4_), .CO(
        u5_mult_82_CARRYB_47__3_), .S(u5_mult_82_SUMB_47__3_) );
  FA_X1 u5_mult_82_S2_47_2 ( .A(u5_mult_82_ab_47__2_), .B(
        u5_mult_82_CARRYB_46__2_), .CI(u5_mult_82_SUMB_46__3_), .CO(
        u5_mult_82_CARRYB_47__2_), .S(u5_mult_82_SUMB_47__2_) );
  FA_X1 u5_mult_82_S2_47_1 ( .A(u5_mult_82_ab_47__1_), .B(
        u5_mult_82_CARRYB_46__1_), .CI(u5_mult_82_SUMB_46__2_), .CO(
        u5_mult_82_CARRYB_47__1_), .S(u5_mult_82_SUMB_47__1_) );
  FA_X1 u5_mult_82_S1_47_0 ( .A(u5_mult_82_ab_47__0_), .B(
        u5_mult_82_CARRYB_46__0_), .CI(u5_mult_82_SUMB_46__1_), .CO(
        u5_mult_82_CARRYB_47__0_), .S(u5_N47) );
  FA_X1 u5_mult_82_S3_48_51 ( .A(u5_mult_82_ab_48__51_), .B(
        u5_mult_82_CARRYB_47__51_), .CI(u5_mult_82_ab_47__52_), .CO(
        u5_mult_82_CARRYB_48__51_), .S(u5_mult_82_SUMB_48__51_) );
  FA_X1 u5_mult_82_S2_48_50 ( .A(u5_mult_82_ab_48__50_), .B(
        u5_mult_82_CARRYB_47__50_), .CI(u5_mult_82_SUMB_47__51_), .CO(
        u5_mult_82_CARRYB_48__50_), .S(u5_mult_82_SUMB_48__50_) );
  FA_X1 u5_mult_82_S2_48_49 ( .A(u5_mult_82_ab_48__49_), .B(
        u5_mult_82_CARRYB_47__49_), .CI(u5_mult_82_SUMB_47__50_), .CO(
        u5_mult_82_CARRYB_48__49_), .S(u5_mult_82_SUMB_48__49_) );
  FA_X1 u5_mult_82_S2_48_48 ( .A(u5_mult_82_ab_48__48_), .B(
        u5_mult_82_CARRYB_47__48_), .CI(u5_mult_82_SUMB_47__49_), .CO(
        u5_mult_82_CARRYB_48__48_), .S(u5_mult_82_SUMB_48__48_) );
  FA_X1 u5_mult_82_S2_48_47 ( .A(u5_mult_82_ab_48__47_), .B(
        u5_mult_82_CARRYB_47__47_), .CI(u5_mult_82_SUMB_47__48_), .CO(
        u5_mult_82_CARRYB_48__47_), .S(u5_mult_82_SUMB_48__47_) );
  FA_X1 u5_mult_82_S2_48_46 ( .A(u5_mult_82_ab_48__46_), .B(
        u5_mult_82_CARRYB_47__46_), .CI(u5_mult_82_SUMB_47__47_), .CO(
        u5_mult_82_CARRYB_48__46_), .S(u5_mult_82_SUMB_48__46_) );
  FA_X1 u5_mult_82_S2_48_45 ( .A(u5_mult_82_ab_48__45_), .B(
        u5_mult_82_CARRYB_47__45_), .CI(u5_mult_82_SUMB_47__46_), .CO(
        u5_mult_82_CARRYB_48__45_), .S(u5_mult_82_SUMB_48__45_) );
  FA_X1 u5_mult_82_S2_48_44 ( .A(u5_mult_82_ab_48__44_), .B(
        u5_mult_82_CARRYB_47__44_), .CI(u5_mult_82_SUMB_47__45_), .CO(
        u5_mult_82_CARRYB_48__44_), .S(u5_mult_82_SUMB_48__44_) );
  FA_X1 u5_mult_82_S2_48_43 ( .A(u5_mult_82_ab_48__43_), .B(
        u5_mult_82_CARRYB_47__43_), .CI(u5_mult_82_SUMB_47__44_), .CO(
        u5_mult_82_CARRYB_48__43_), .S(u5_mult_82_SUMB_48__43_) );
  FA_X1 u5_mult_82_S2_48_42 ( .A(u5_mult_82_ab_48__42_), .B(
        u5_mult_82_CARRYB_47__42_), .CI(u5_mult_82_SUMB_47__43_), .CO(
        u5_mult_82_CARRYB_48__42_), .S(u5_mult_82_SUMB_48__42_) );
  FA_X1 u5_mult_82_S2_48_41 ( .A(u5_mult_82_ab_48__41_), .B(
        u5_mult_82_CARRYB_47__41_), .CI(u5_mult_82_SUMB_47__42_), .CO(
        u5_mult_82_CARRYB_48__41_), .S(u5_mult_82_SUMB_48__41_) );
  FA_X1 u5_mult_82_S2_48_40 ( .A(u5_mult_82_ab_48__40_), .B(
        u5_mult_82_CARRYB_47__40_), .CI(u5_mult_82_SUMB_47__41_), .CO(
        u5_mult_82_CARRYB_48__40_), .S(u5_mult_82_SUMB_48__40_) );
  FA_X1 u5_mult_82_S2_48_39 ( .A(u5_mult_82_ab_48__39_), .B(
        u5_mult_82_CARRYB_47__39_), .CI(u5_mult_82_SUMB_47__40_), .CO(
        u5_mult_82_CARRYB_48__39_), .S(u5_mult_82_SUMB_48__39_) );
  FA_X1 u5_mult_82_S2_48_38 ( .A(u5_mult_82_ab_48__38_), .B(
        u5_mult_82_CARRYB_47__38_), .CI(u5_mult_82_SUMB_47__39_), .CO(
        u5_mult_82_CARRYB_48__38_), .S(u5_mult_82_SUMB_48__38_) );
  FA_X1 u5_mult_82_S2_48_37 ( .A(u5_mult_82_ab_48__37_), .B(
        u5_mult_82_CARRYB_47__37_), .CI(u5_mult_82_SUMB_47__38_), .CO(
        u5_mult_82_CARRYB_48__37_), .S(u5_mult_82_SUMB_48__37_) );
  FA_X1 u5_mult_82_S2_48_36 ( .A(u5_mult_82_ab_48__36_), .B(
        u5_mult_82_CARRYB_47__36_), .CI(u5_mult_82_SUMB_47__37_), .CO(
        u5_mult_82_CARRYB_48__36_), .S(u5_mult_82_SUMB_48__36_) );
  FA_X1 u5_mult_82_S2_48_35 ( .A(u5_mult_82_ab_48__35_), .B(
        u5_mult_82_CARRYB_47__35_), .CI(u5_mult_82_SUMB_47__36_), .CO(
        u5_mult_82_CARRYB_48__35_), .S(u5_mult_82_SUMB_48__35_) );
  FA_X1 u5_mult_82_S2_48_34 ( .A(u5_mult_82_ab_48__34_), .B(
        u5_mult_82_CARRYB_47__34_), .CI(u5_mult_82_SUMB_47__35_), .CO(
        u5_mult_82_CARRYB_48__34_), .S(u5_mult_82_SUMB_48__34_) );
  FA_X1 u5_mult_82_S2_48_33 ( .A(u5_mult_82_ab_48__33_), .B(
        u5_mult_82_CARRYB_47__33_), .CI(u5_mult_82_SUMB_47__34_), .CO(
        u5_mult_82_CARRYB_48__33_), .S(u5_mult_82_SUMB_48__33_) );
  FA_X1 u5_mult_82_S2_48_32 ( .A(u5_mult_82_ab_48__32_), .B(
        u5_mult_82_CARRYB_47__32_), .CI(u5_mult_82_SUMB_47__33_), .CO(
        u5_mult_82_CARRYB_48__32_), .S(u5_mult_82_SUMB_48__32_) );
  FA_X1 u5_mult_82_S2_48_31 ( .A(u5_mult_82_ab_48__31_), .B(
        u5_mult_82_CARRYB_47__31_), .CI(u5_mult_82_SUMB_47__32_), .CO(
        u5_mult_82_CARRYB_48__31_), .S(u5_mult_82_SUMB_48__31_) );
  FA_X1 u5_mult_82_S2_48_30 ( .A(u5_mult_82_ab_48__30_), .B(
        u5_mult_82_CARRYB_47__30_), .CI(u5_mult_82_SUMB_47__31_), .CO(
        u5_mult_82_CARRYB_48__30_), .S(u5_mult_82_SUMB_48__30_) );
  FA_X1 u5_mult_82_S2_48_29 ( .A(u5_mult_82_ab_48__29_), .B(
        u5_mult_82_CARRYB_47__29_), .CI(u5_mult_82_SUMB_47__30_), .CO(
        u5_mult_82_CARRYB_48__29_), .S(u5_mult_82_SUMB_48__29_) );
  FA_X1 u5_mult_82_S2_48_28 ( .A(u5_mult_82_ab_48__28_), .B(
        u5_mult_82_CARRYB_47__28_), .CI(u5_mult_82_SUMB_47__29_), .CO(
        u5_mult_82_CARRYB_48__28_), .S(u5_mult_82_SUMB_48__28_) );
  FA_X1 u5_mult_82_S2_48_27 ( .A(u5_mult_82_ab_48__27_), .B(
        u5_mult_82_CARRYB_47__27_), .CI(u5_mult_82_SUMB_47__28_), .CO(
        u5_mult_82_CARRYB_48__27_), .S(u5_mult_82_SUMB_48__27_) );
  FA_X1 u5_mult_82_S2_48_26 ( .A(u5_mult_82_ab_48__26_), .B(
        u5_mult_82_CARRYB_47__26_), .CI(u5_mult_82_SUMB_47__27_), .CO(
        u5_mult_82_CARRYB_48__26_), .S(u5_mult_82_SUMB_48__26_) );
  FA_X1 u5_mult_82_S2_48_25 ( .A(u5_mult_82_ab_48__25_), .B(
        u5_mult_82_CARRYB_47__25_), .CI(u5_mult_82_SUMB_47__26_), .CO(
        u5_mult_82_CARRYB_48__25_), .S(u5_mult_82_SUMB_48__25_) );
  FA_X1 u5_mult_82_S2_48_24 ( .A(u5_mult_82_ab_48__24_), .B(
        u5_mult_82_CARRYB_47__24_), .CI(u5_mult_82_SUMB_47__25_), .CO(
        u5_mult_82_CARRYB_48__24_), .S(u5_mult_82_SUMB_48__24_) );
  FA_X1 u5_mult_82_S2_48_23 ( .A(u5_mult_82_ab_48__23_), .B(
        u5_mult_82_CARRYB_47__23_), .CI(u5_mult_82_SUMB_47__24_), .CO(
        u5_mult_82_CARRYB_48__23_), .S(u5_mult_82_SUMB_48__23_) );
  FA_X1 u5_mult_82_S2_48_22 ( .A(u5_mult_82_ab_48__22_), .B(
        u5_mult_82_CARRYB_47__22_), .CI(u5_mult_82_SUMB_47__23_), .CO(
        u5_mult_82_CARRYB_48__22_), .S(u5_mult_82_SUMB_48__22_) );
  FA_X1 u5_mult_82_S2_48_21 ( .A(u5_mult_82_ab_48__21_), .B(
        u5_mult_82_CARRYB_47__21_), .CI(u5_mult_82_SUMB_47__22_), .CO(
        u5_mult_82_CARRYB_48__21_), .S(u5_mult_82_SUMB_48__21_) );
  FA_X1 u5_mult_82_S2_48_20 ( .A(u5_mult_82_ab_48__20_), .B(
        u5_mult_82_CARRYB_47__20_), .CI(u5_mult_82_SUMB_47__21_), .CO(
        u5_mult_82_CARRYB_48__20_), .S(u5_mult_82_SUMB_48__20_) );
  FA_X1 u5_mult_82_S2_48_19 ( .A(u5_mult_82_ab_48__19_), .B(
        u5_mult_82_CARRYB_47__19_), .CI(u5_mult_82_SUMB_47__20_), .CO(
        u5_mult_82_CARRYB_48__19_), .S(u5_mult_82_SUMB_48__19_) );
  FA_X1 u5_mult_82_S2_48_18 ( .A(u5_mult_82_ab_48__18_), .B(
        u5_mult_82_CARRYB_47__18_), .CI(u5_mult_82_SUMB_47__19_), .CO(
        u5_mult_82_CARRYB_48__18_), .S(u5_mult_82_SUMB_48__18_) );
  FA_X1 u5_mult_82_S2_48_17 ( .A(u5_mult_82_ab_48__17_), .B(
        u5_mult_82_CARRYB_47__17_), .CI(u5_mult_82_SUMB_47__18_), .CO(
        u5_mult_82_CARRYB_48__17_), .S(u5_mult_82_SUMB_48__17_) );
  FA_X1 u5_mult_82_S2_48_16 ( .A(u5_mult_82_ab_48__16_), .B(
        u5_mult_82_CARRYB_47__16_), .CI(u5_mult_82_SUMB_47__17_), .CO(
        u5_mult_82_CARRYB_48__16_), .S(u5_mult_82_SUMB_48__16_) );
  FA_X1 u5_mult_82_S2_48_15 ( .A(u5_mult_82_ab_48__15_), .B(
        u5_mult_82_CARRYB_47__15_), .CI(u5_mult_82_SUMB_47__16_), .CO(
        u5_mult_82_CARRYB_48__15_), .S(u5_mult_82_SUMB_48__15_) );
  FA_X1 u5_mult_82_S2_48_14 ( .A(u5_mult_82_ab_48__14_), .B(
        u5_mult_82_CARRYB_47__14_), .CI(u5_mult_82_SUMB_47__15_), .CO(
        u5_mult_82_CARRYB_48__14_), .S(u5_mult_82_SUMB_48__14_) );
  FA_X1 u5_mult_82_S2_48_13 ( .A(u5_mult_82_ab_48__13_), .B(
        u5_mult_82_CARRYB_47__13_), .CI(u5_mult_82_SUMB_47__14_), .CO(
        u5_mult_82_CARRYB_48__13_), .S(u5_mult_82_SUMB_48__13_) );
  FA_X1 u5_mult_82_S2_48_12 ( .A(u5_mult_82_ab_48__12_), .B(
        u5_mult_82_CARRYB_47__12_), .CI(u5_mult_82_SUMB_47__13_), .CO(
        u5_mult_82_CARRYB_48__12_), .S(u5_mult_82_SUMB_48__12_) );
  FA_X1 u5_mult_82_S2_48_11 ( .A(u5_mult_82_ab_48__11_), .B(
        u5_mult_82_CARRYB_47__11_), .CI(u5_mult_82_SUMB_47__12_), .CO(
        u5_mult_82_CARRYB_48__11_), .S(u5_mult_82_SUMB_48__11_) );
  FA_X1 u5_mult_82_S2_48_10 ( .A(u5_mult_82_ab_48__10_), .B(
        u5_mult_82_CARRYB_47__10_), .CI(u5_mult_82_SUMB_47__11_), .CO(
        u5_mult_82_CARRYB_48__10_), .S(u5_mult_82_SUMB_48__10_) );
  FA_X1 u5_mult_82_S2_48_9 ( .A(u5_mult_82_ab_48__9_), .B(
        u5_mult_82_CARRYB_47__9_), .CI(u5_mult_82_SUMB_47__10_), .CO(
        u5_mult_82_CARRYB_48__9_), .S(u5_mult_82_SUMB_48__9_) );
  FA_X1 u5_mult_82_S2_48_8 ( .A(u5_mult_82_ab_48__8_), .B(
        u5_mult_82_CARRYB_47__8_), .CI(u5_mult_82_SUMB_47__9_), .CO(
        u5_mult_82_CARRYB_48__8_), .S(u5_mult_82_SUMB_48__8_) );
  FA_X1 u5_mult_82_S2_48_7 ( .A(u5_mult_82_ab_48__7_), .B(
        u5_mult_82_CARRYB_47__7_), .CI(u5_mult_82_SUMB_47__8_), .CO(
        u5_mult_82_CARRYB_48__7_), .S(u5_mult_82_SUMB_48__7_) );
  FA_X1 u5_mult_82_S2_48_6 ( .A(u5_mult_82_ab_48__6_), .B(
        u5_mult_82_CARRYB_47__6_), .CI(u5_mult_82_SUMB_47__7_), .CO(
        u5_mult_82_CARRYB_48__6_), .S(u5_mult_82_SUMB_48__6_) );
  FA_X1 u5_mult_82_S2_48_5 ( .A(u5_mult_82_ab_48__5_), .B(
        u5_mult_82_CARRYB_47__5_), .CI(u5_mult_82_SUMB_47__6_), .CO(
        u5_mult_82_CARRYB_48__5_), .S(u5_mult_82_SUMB_48__5_) );
  FA_X1 u5_mult_82_S2_48_4 ( .A(u5_mult_82_ab_48__4_), .B(
        u5_mult_82_CARRYB_47__4_), .CI(u5_mult_82_SUMB_47__5_), .CO(
        u5_mult_82_CARRYB_48__4_), .S(u5_mult_82_SUMB_48__4_) );
  FA_X1 u5_mult_82_S2_48_3 ( .A(u5_mult_82_ab_48__3_), .B(
        u5_mult_82_CARRYB_47__3_), .CI(u5_mult_82_SUMB_47__4_), .CO(
        u5_mult_82_CARRYB_48__3_), .S(u5_mult_82_SUMB_48__3_) );
  FA_X1 u5_mult_82_S2_48_2 ( .A(u5_mult_82_ab_48__2_), .B(
        u5_mult_82_CARRYB_47__2_), .CI(u5_mult_82_SUMB_47__3_), .CO(
        u5_mult_82_CARRYB_48__2_), .S(u5_mult_82_SUMB_48__2_) );
  FA_X1 u5_mult_82_S2_48_1 ( .A(u5_mult_82_ab_48__1_), .B(
        u5_mult_82_CARRYB_47__1_), .CI(u5_mult_82_SUMB_47__2_), .CO(
        u5_mult_82_CARRYB_48__1_), .S(u5_mult_82_SUMB_48__1_) );
  FA_X1 u5_mult_82_S1_48_0 ( .A(u5_mult_82_ab_48__0_), .B(
        u5_mult_82_CARRYB_47__0_), .CI(u5_mult_82_SUMB_47__1_), .CO(
        u5_mult_82_CARRYB_48__0_), .S(u5_N48) );
  FA_X1 u5_mult_82_S3_49_51 ( .A(u5_mult_82_ab_49__51_), .B(
        u5_mult_82_CARRYB_48__51_), .CI(u5_mult_82_ab_48__52_), .CO(
        u5_mult_82_CARRYB_49__51_), .S(u5_mult_82_SUMB_49__51_) );
  FA_X1 u5_mult_82_S2_49_50 ( .A(u5_mult_82_ab_49__50_), .B(
        u5_mult_82_CARRYB_48__50_), .CI(u5_mult_82_SUMB_48__51_), .CO(
        u5_mult_82_CARRYB_49__50_), .S(u5_mult_82_SUMB_49__50_) );
  FA_X1 u5_mult_82_S2_49_49 ( .A(u5_mult_82_ab_49__49_), .B(
        u5_mult_82_CARRYB_48__49_), .CI(u5_mult_82_SUMB_48__50_), .CO(
        u5_mult_82_CARRYB_49__49_), .S(u5_mult_82_SUMB_49__49_) );
  FA_X1 u5_mult_82_S2_49_48 ( .A(u5_mult_82_ab_49__48_), .B(
        u5_mult_82_CARRYB_48__48_), .CI(u5_mult_82_SUMB_48__49_), .CO(
        u5_mult_82_CARRYB_49__48_), .S(u5_mult_82_SUMB_49__48_) );
  FA_X1 u5_mult_82_S2_49_47 ( .A(u5_mult_82_ab_49__47_), .B(
        u5_mult_82_CARRYB_48__47_), .CI(u5_mult_82_SUMB_48__48_), .CO(
        u5_mult_82_CARRYB_49__47_), .S(u5_mult_82_SUMB_49__47_) );
  FA_X1 u5_mult_82_S2_49_46 ( .A(u5_mult_82_ab_49__46_), .B(
        u5_mult_82_CARRYB_48__46_), .CI(u5_mult_82_SUMB_48__47_), .CO(
        u5_mult_82_CARRYB_49__46_), .S(u5_mult_82_SUMB_49__46_) );
  FA_X1 u5_mult_82_S2_49_45 ( .A(u5_mult_82_ab_49__45_), .B(
        u5_mult_82_CARRYB_48__45_), .CI(u5_mult_82_SUMB_48__46_), .CO(
        u5_mult_82_CARRYB_49__45_), .S(u5_mult_82_SUMB_49__45_) );
  FA_X1 u5_mult_82_S2_49_44 ( .A(u5_mult_82_ab_49__44_), .B(
        u5_mult_82_CARRYB_48__44_), .CI(u5_mult_82_SUMB_48__45_), .CO(
        u5_mult_82_CARRYB_49__44_), .S(u5_mult_82_SUMB_49__44_) );
  FA_X1 u5_mult_82_S2_49_43 ( .A(u5_mult_82_ab_49__43_), .B(
        u5_mult_82_CARRYB_48__43_), .CI(u5_mult_82_SUMB_48__44_), .CO(
        u5_mult_82_CARRYB_49__43_), .S(u5_mult_82_SUMB_49__43_) );
  FA_X1 u5_mult_82_S2_49_42 ( .A(u5_mult_82_ab_49__42_), .B(
        u5_mult_82_CARRYB_48__42_), .CI(u5_mult_82_SUMB_48__43_), .CO(
        u5_mult_82_CARRYB_49__42_), .S(u5_mult_82_SUMB_49__42_) );
  FA_X1 u5_mult_82_S2_49_41 ( .A(u5_mult_82_ab_49__41_), .B(
        u5_mult_82_CARRYB_48__41_), .CI(u5_mult_82_SUMB_48__42_), .CO(
        u5_mult_82_CARRYB_49__41_), .S(u5_mult_82_SUMB_49__41_) );
  FA_X1 u5_mult_82_S2_49_40 ( .A(u5_mult_82_ab_49__40_), .B(
        u5_mult_82_CARRYB_48__40_), .CI(u5_mult_82_SUMB_48__41_), .CO(
        u5_mult_82_CARRYB_49__40_), .S(u5_mult_82_SUMB_49__40_) );
  FA_X1 u5_mult_82_S2_49_39 ( .A(u5_mult_82_ab_49__39_), .B(
        u5_mult_82_CARRYB_48__39_), .CI(u5_mult_82_SUMB_48__40_), .CO(
        u5_mult_82_CARRYB_49__39_), .S(u5_mult_82_SUMB_49__39_) );
  FA_X1 u5_mult_82_S2_49_38 ( .A(u5_mult_82_ab_49__38_), .B(
        u5_mult_82_CARRYB_48__38_), .CI(u5_mult_82_SUMB_48__39_), .CO(
        u5_mult_82_CARRYB_49__38_), .S(u5_mult_82_SUMB_49__38_) );
  FA_X1 u5_mult_82_S2_49_37 ( .A(u5_mult_82_ab_49__37_), .B(
        u5_mult_82_CARRYB_48__37_), .CI(u5_mult_82_SUMB_48__38_), .CO(
        u5_mult_82_CARRYB_49__37_), .S(u5_mult_82_SUMB_49__37_) );
  FA_X1 u5_mult_82_S2_49_36 ( .A(u5_mult_82_ab_49__36_), .B(
        u5_mult_82_CARRYB_48__36_), .CI(u5_mult_82_SUMB_48__37_), .CO(
        u5_mult_82_CARRYB_49__36_), .S(u5_mult_82_SUMB_49__36_) );
  FA_X1 u5_mult_82_S2_49_35 ( .A(u5_mult_82_ab_49__35_), .B(
        u5_mult_82_CARRYB_48__35_), .CI(u5_mult_82_SUMB_48__36_), .CO(
        u5_mult_82_CARRYB_49__35_), .S(u5_mult_82_SUMB_49__35_) );
  FA_X1 u5_mult_82_S2_49_34 ( .A(u5_mult_82_ab_49__34_), .B(
        u5_mult_82_CARRYB_48__34_), .CI(u5_mult_82_SUMB_48__35_), .CO(
        u5_mult_82_CARRYB_49__34_), .S(u5_mult_82_SUMB_49__34_) );
  FA_X1 u5_mult_82_S2_49_33 ( .A(u5_mult_82_ab_49__33_), .B(
        u5_mult_82_CARRYB_48__33_), .CI(u5_mult_82_SUMB_48__34_), .CO(
        u5_mult_82_CARRYB_49__33_), .S(u5_mult_82_SUMB_49__33_) );
  FA_X1 u5_mult_82_S2_49_32 ( .A(u5_mult_82_ab_49__32_), .B(
        u5_mult_82_CARRYB_48__32_), .CI(u5_mult_82_SUMB_48__33_), .CO(
        u5_mult_82_CARRYB_49__32_), .S(u5_mult_82_SUMB_49__32_) );
  FA_X1 u5_mult_82_S2_49_31 ( .A(u5_mult_82_ab_49__31_), .B(
        u5_mult_82_CARRYB_48__31_), .CI(u5_mult_82_SUMB_48__32_), .CO(
        u5_mult_82_CARRYB_49__31_), .S(u5_mult_82_SUMB_49__31_) );
  FA_X1 u5_mult_82_S2_49_30 ( .A(u5_mult_82_ab_49__30_), .B(
        u5_mult_82_CARRYB_48__30_), .CI(u5_mult_82_SUMB_48__31_), .CO(
        u5_mult_82_CARRYB_49__30_), .S(u5_mult_82_SUMB_49__30_) );
  FA_X1 u5_mult_82_S2_49_29 ( .A(u5_mult_82_ab_49__29_), .B(
        u5_mult_82_CARRYB_48__29_), .CI(u5_mult_82_SUMB_48__30_), .CO(
        u5_mult_82_CARRYB_49__29_), .S(u5_mult_82_SUMB_49__29_) );
  FA_X1 u5_mult_82_S2_49_28 ( .A(u5_mult_82_ab_49__28_), .B(
        u5_mult_82_CARRYB_48__28_), .CI(u5_mult_82_SUMB_48__29_), .CO(
        u5_mult_82_CARRYB_49__28_), .S(u5_mult_82_SUMB_49__28_) );
  FA_X1 u5_mult_82_S2_49_27 ( .A(u5_mult_82_ab_49__27_), .B(
        u5_mult_82_CARRYB_48__27_), .CI(u5_mult_82_SUMB_48__28_), .CO(
        u5_mult_82_CARRYB_49__27_), .S(u5_mult_82_SUMB_49__27_) );
  FA_X1 u5_mult_82_S2_49_26 ( .A(u5_mult_82_ab_49__26_), .B(
        u5_mult_82_CARRYB_48__26_), .CI(u5_mult_82_SUMB_48__27_), .CO(
        u5_mult_82_CARRYB_49__26_), .S(u5_mult_82_SUMB_49__26_) );
  FA_X1 u5_mult_82_S2_49_25 ( .A(u5_mult_82_ab_49__25_), .B(
        u5_mult_82_CARRYB_48__25_), .CI(u5_mult_82_SUMB_48__26_), .CO(
        u5_mult_82_CARRYB_49__25_), .S(u5_mult_82_SUMB_49__25_) );
  FA_X1 u5_mult_82_S2_49_24 ( .A(u5_mult_82_ab_49__24_), .B(
        u5_mult_82_CARRYB_48__24_), .CI(u5_mult_82_SUMB_48__25_), .CO(
        u5_mult_82_CARRYB_49__24_), .S(u5_mult_82_SUMB_49__24_) );
  FA_X1 u5_mult_82_S2_49_23 ( .A(u5_mult_82_ab_49__23_), .B(
        u5_mult_82_CARRYB_48__23_), .CI(u5_mult_82_SUMB_48__24_), .CO(
        u5_mult_82_CARRYB_49__23_), .S(u5_mult_82_SUMB_49__23_) );
  FA_X1 u5_mult_82_S2_49_22 ( .A(u5_mult_82_ab_49__22_), .B(
        u5_mult_82_CARRYB_48__22_), .CI(u5_mult_82_SUMB_48__23_), .CO(
        u5_mult_82_CARRYB_49__22_), .S(u5_mult_82_SUMB_49__22_) );
  FA_X1 u5_mult_82_S2_49_21 ( .A(u5_mult_82_ab_49__21_), .B(
        u5_mult_82_CARRYB_48__21_), .CI(u5_mult_82_SUMB_48__22_), .CO(
        u5_mult_82_CARRYB_49__21_), .S(u5_mult_82_SUMB_49__21_) );
  FA_X1 u5_mult_82_S2_49_20 ( .A(u5_mult_82_ab_49__20_), .B(
        u5_mult_82_CARRYB_48__20_), .CI(u5_mult_82_SUMB_48__21_), .CO(
        u5_mult_82_CARRYB_49__20_), .S(u5_mult_82_SUMB_49__20_) );
  FA_X1 u5_mult_82_S2_49_19 ( .A(u5_mult_82_ab_49__19_), .B(
        u5_mult_82_CARRYB_48__19_), .CI(u5_mult_82_SUMB_48__20_), .CO(
        u5_mult_82_CARRYB_49__19_), .S(u5_mult_82_SUMB_49__19_) );
  FA_X1 u5_mult_82_S2_49_18 ( .A(u5_mult_82_ab_49__18_), .B(
        u5_mult_82_CARRYB_48__18_), .CI(u5_mult_82_SUMB_48__19_), .CO(
        u5_mult_82_CARRYB_49__18_), .S(u5_mult_82_SUMB_49__18_) );
  FA_X1 u5_mult_82_S2_49_17 ( .A(u5_mult_82_ab_49__17_), .B(
        u5_mult_82_CARRYB_48__17_), .CI(u5_mult_82_SUMB_48__18_), .CO(
        u5_mult_82_CARRYB_49__17_), .S(u5_mult_82_SUMB_49__17_) );
  FA_X1 u5_mult_82_S2_49_16 ( .A(u5_mult_82_ab_49__16_), .B(
        u5_mult_82_CARRYB_48__16_), .CI(u5_mult_82_SUMB_48__17_), .CO(
        u5_mult_82_CARRYB_49__16_), .S(u5_mult_82_SUMB_49__16_) );
  FA_X1 u5_mult_82_S2_49_15 ( .A(u5_mult_82_ab_49__15_), .B(
        u5_mult_82_CARRYB_48__15_), .CI(u5_mult_82_SUMB_48__16_), .CO(
        u5_mult_82_CARRYB_49__15_), .S(u5_mult_82_SUMB_49__15_) );
  FA_X1 u5_mult_82_S2_49_14 ( .A(u5_mult_82_ab_49__14_), .B(
        u5_mult_82_CARRYB_48__14_), .CI(u5_mult_82_SUMB_48__15_), .CO(
        u5_mult_82_CARRYB_49__14_), .S(u5_mult_82_SUMB_49__14_) );
  FA_X1 u5_mult_82_S2_49_13 ( .A(u5_mult_82_ab_49__13_), .B(
        u5_mult_82_CARRYB_48__13_), .CI(u5_mult_82_SUMB_48__14_), .CO(
        u5_mult_82_CARRYB_49__13_), .S(u5_mult_82_SUMB_49__13_) );
  FA_X1 u5_mult_82_S2_49_12 ( .A(u5_mult_82_ab_49__12_), .B(
        u5_mult_82_CARRYB_48__12_), .CI(u5_mult_82_SUMB_48__13_), .CO(
        u5_mult_82_CARRYB_49__12_), .S(u5_mult_82_SUMB_49__12_) );
  FA_X1 u5_mult_82_S2_49_11 ( .A(u5_mult_82_ab_49__11_), .B(
        u5_mult_82_CARRYB_48__11_), .CI(u5_mult_82_SUMB_48__12_), .CO(
        u5_mult_82_CARRYB_49__11_), .S(u5_mult_82_SUMB_49__11_) );
  FA_X1 u5_mult_82_S2_49_10 ( .A(u5_mult_82_ab_49__10_), .B(
        u5_mult_82_CARRYB_48__10_), .CI(u5_mult_82_SUMB_48__11_), .CO(
        u5_mult_82_CARRYB_49__10_), .S(u5_mult_82_SUMB_49__10_) );
  FA_X1 u5_mult_82_S2_49_9 ( .A(u5_mult_82_ab_49__9_), .B(
        u5_mult_82_CARRYB_48__9_), .CI(u5_mult_82_SUMB_48__10_), .CO(
        u5_mult_82_CARRYB_49__9_), .S(u5_mult_82_SUMB_49__9_) );
  FA_X1 u5_mult_82_S2_49_8 ( .A(u5_mult_82_ab_49__8_), .B(
        u5_mult_82_CARRYB_48__8_), .CI(u5_mult_82_SUMB_48__9_), .CO(
        u5_mult_82_CARRYB_49__8_), .S(u5_mult_82_SUMB_49__8_) );
  FA_X1 u5_mult_82_S2_49_7 ( .A(u5_mult_82_ab_49__7_), .B(
        u5_mult_82_CARRYB_48__7_), .CI(u5_mult_82_SUMB_48__8_), .CO(
        u5_mult_82_CARRYB_49__7_), .S(u5_mult_82_SUMB_49__7_) );
  FA_X1 u5_mult_82_S2_49_6 ( .A(u5_mult_82_ab_49__6_), .B(
        u5_mult_82_CARRYB_48__6_), .CI(u5_mult_82_SUMB_48__7_), .CO(
        u5_mult_82_CARRYB_49__6_), .S(u5_mult_82_SUMB_49__6_) );
  FA_X1 u5_mult_82_S2_49_5 ( .A(u5_mult_82_ab_49__5_), .B(
        u5_mult_82_CARRYB_48__5_), .CI(u5_mult_82_SUMB_48__6_), .CO(
        u5_mult_82_CARRYB_49__5_), .S(u5_mult_82_SUMB_49__5_) );
  FA_X1 u5_mult_82_S2_49_4 ( .A(u5_mult_82_ab_49__4_), .B(
        u5_mult_82_CARRYB_48__4_), .CI(u5_mult_82_SUMB_48__5_), .CO(
        u5_mult_82_CARRYB_49__4_), .S(u5_mult_82_SUMB_49__4_) );
  FA_X1 u5_mult_82_S2_49_3 ( .A(u5_mult_82_ab_49__3_), .B(
        u5_mult_82_CARRYB_48__3_), .CI(u5_mult_82_SUMB_48__4_), .CO(
        u5_mult_82_CARRYB_49__3_), .S(u5_mult_82_SUMB_49__3_) );
  FA_X1 u5_mult_82_S2_49_2 ( .A(u5_mult_82_ab_49__2_), .B(
        u5_mult_82_CARRYB_48__2_), .CI(u5_mult_82_SUMB_48__3_), .CO(
        u5_mult_82_CARRYB_49__2_), .S(u5_mult_82_SUMB_49__2_) );
  FA_X1 u5_mult_82_S2_49_1 ( .A(u5_mult_82_ab_49__1_), .B(
        u5_mult_82_CARRYB_48__1_), .CI(u5_mult_82_SUMB_48__2_), .CO(
        u5_mult_82_CARRYB_49__1_), .S(u5_mult_82_SUMB_49__1_) );
  FA_X1 u5_mult_82_S1_49_0 ( .A(u5_mult_82_ab_49__0_), .B(
        u5_mult_82_CARRYB_48__0_), .CI(u5_mult_82_SUMB_48__1_), .CO(
        u5_mult_82_CARRYB_49__0_), .S(u5_N49) );
  FA_X1 u5_mult_82_S3_50_51 ( .A(u5_mult_82_ab_50__51_), .B(
        u5_mult_82_CARRYB_49__51_), .CI(u5_mult_82_ab_49__52_), .CO(
        u5_mult_82_CARRYB_50__51_), .S(u5_mult_82_SUMB_50__51_) );
  FA_X1 u5_mult_82_S2_50_50 ( .A(u5_mult_82_ab_50__50_), .B(
        u5_mult_82_CARRYB_49__50_), .CI(u5_mult_82_SUMB_49__51_), .CO(
        u5_mult_82_CARRYB_50__50_), .S(u5_mult_82_SUMB_50__50_) );
  FA_X1 u5_mult_82_S2_50_49 ( .A(u5_mult_82_ab_50__49_), .B(
        u5_mult_82_CARRYB_49__49_), .CI(u5_mult_82_SUMB_49__50_), .CO(
        u5_mult_82_CARRYB_50__49_), .S(u5_mult_82_SUMB_50__49_) );
  FA_X1 u5_mult_82_S2_50_48 ( .A(u5_mult_82_ab_50__48_), .B(
        u5_mult_82_CARRYB_49__48_), .CI(u5_mult_82_SUMB_49__49_), .CO(
        u5_mult_82_CARRYB_50__48_), .S(u5_mult_82_SUMB_50__48_) );
  FA_X1 u5_mult_82_S2_50_47 ( .A(u5_mult_82_ab_50__47_), .B(
        u5_mult_82_CARRYB_49__47_), .CI(u5_mult_82_SUMB_49__48_), .CO(
        u5_mult_82_CARRYB_50__47_), .S(u5_mult_82_SUMB_50__47_) );
  FA_X1 u5_mult_82_S2_50_46 ( .A(u5_mult_82_ab_50__46_), .B(
        u5_mult_82_CARRYB_49__46_), .CI(u5_mult_82_SUMB_49__47_), .CO(
        u5_mult_82_CARRYB_50__46_), .S(u5_mult_82_SUMB_50__46_) );
  FA_X1 u5_mult_82_S2_50_45 ( .A(u5_mult_82_ab_50__45_), .B(
        u5_mult_82_CARRYB_49__45_), .CI(u5_mult_82_SUMB_49__46_), .CO(
        u5_mult_82_CARRYB_50__45_), .S(u5_mult_82_SUMB_50__45_) );
  FA_X1 u5_mult_82_S2_50_44 ( .A(u5_mult_82_ab_50__44_), .B(
        u5_mult_82_CARRYB_49__44_), .CI(u5_mult_82_SUMB_49__45_), .CO(
        u5_mult_82_CARRYB_50__44_), .S(u5_mult_82_SUMB_50__44_) );
  FA_X1 u5_mult_82_S2_50_43 ( .A(u5_mult_82_ab_50__43_), .B(
        u5_mult_82_CARRYB_49__43_), .CI(u5_mult_82_SUMB_49__44_), .CO(
        u5_mult_82_CARRYB_50__43_), .S(u5_mult_82_SUMB_50__43_) );
  FA_X1 u5_mult_82_S2_50_42 ( .A(u5_mult_82_ab_50__42_), .B(
        u5_mult_82_CARRYB_49__42_), .CI(u5_mult_82_SUMB_49__43_), .CO(
        u5_mult_82_CARRYB_50__42_), .S(u5_mult_82_SUMB_50__42_) );
  FA_X1 u5_mult_82_S2_50_41 ( .A(u5_mult_82_ab_50__41_), .B(
        u5_mult_82_CARRYB_49__41_), .CI(u5_mult_82_SUMB_49__42_), .CO(
        u5_mult_82_CARRYB_50__41_), .S(u5_mult_82_SUMB_50__41_) );
  FA_X1 u5_mult_82_S2_50_40 ( .A(u5_mult_82_ab_50__40_), .B(
        u5_mult_82_CARRYB_49__40_), .CI(u5_mult_82_SUMB_49__41_), .CO(
        u5_mult_82_CARRYB_50__40_), .S(u5_mult_82_SUMB_50__40_) );
  FA_X1 u5_mult_82_S2_50_39 ( .A(u5_mult_82_ab_50__39_), .B(
        u5_mult_82_CARRYB_49__39_), .CI(u5_mult_82_SUMB_49__40_), .CO(
        u5_mult_82_CARRYB_50__39_), .S(u5_mult_82_SUMB_50__39_) );
  FA_X1 u5_mult_82_S2_50_38 ( .A(u5_mult_82_ab_50__38_), .B(
        u5_mult_82_CARRYB_49__38_), .CI(u5_mult_82_SUMB_49__39_), .CO(
        u5_mult_82_CARRYB_50__38_), .S(u5_mult_82_SUMB_50__38_) );
  FA_X1 u5_mult_82_S2_50_37 ( .A(u5_mult_82_ab_50__37_), .B(
        u5_mult_82_CARRYB_49__37_), .CI(u5_mult_82_SUMB_49__38_), .CO(
        u5_mult_82_CARRYB_50__37_), .S(u5_mult_82_SUMB_50__37_) );
  FA_X1 u5_mult_82_S2_50_36 ( .A(u5_mult_82_ab_50__36_), .B(
        u5_mult_82_CARRYB_49__36_), .CI(u5_mult_82_SUMB_49__37_), .CO(
        u5_mult_82_CARRYB_50__36_), .S(u5_mult_82_SUMB_50__36_) );
  FA_X1 u5_mult_82_S2_50_35 ( .A(u5_mult_82_ab_50__35_), .B(
        u5_mult_82_CARRYB_49__35_), .CI(u5_mult_82_SUMB_49__36_), .CO(
        u5_mult_82_CARRYB_50__35_), .S(u5_mult_82_SUMB_50__35_) );
  FA_X1 u5_mult_82_S2_50_34 ( .A(u5_mult_82_ab_50__34_), .B(
        u5_mult_82_CARRYB_49__34_), .CI(u5_mult_82_SUMB_49__35_), .CO(
        u5_mult_82_CARRYB_50__34_), .S(u5_mult_82_SUMB_50__34_) );
  FA_X1 u5_mult_82_S2_50_33 ( .A(u5_mult_82_ab_50__33_), .B(
        u5_mult_82_CARRYB_49__33_), .CI(u5_mult_82_SUMB_49__34_), .CO(
        u5_mult_82_CARRYB_50__33_), .S(u5_mult_82_SUMB_50__33_) );
  FA_X1 u5_mult_82_S2_50_32 ( .A(u5_mult_82_ab_50__32_), .B(
        u5_mult_82_CARRYB_49__32_), .CI(u5_mult_82_SUMB_49__33_), .CO(
        u5_mult_82_CARRYB_50__32_), .S(u5_mult_82_SUMB_50__32_) );
  FA_X1 u5_mult_82_S2_50_31 ( .A(u5_mult_82_ab_50__31_), .B(
        u5_mult_82_CARRYB_49__31_), .CI(u5_mult_82_SUMB_49__32_), .CO(
        u5_mult_82_CARRYB_50__31_), .S(u5_mult_82_SUMB_50__31_) );
  FA_X1 u5_mult_82_S2_50_30 ( .A(u5_mult_82_ab_50__30_), .B(
        u5_mult_82_CARRYB_49__30_), .CI(u5_mult_82_SUMB_49__31_), .CO(
        u5_mult_82_CARRYB_50__30_), .S(u5_mult_82_SUMB_50__30_) );
  FA_X1 u5_mult_82_S2_50_29 ( .A(u5_mult_82_ab_50__29_), .B(
        u5_mult_82_CARRYB_49__29_), .CI(u5_mult_82_SUMB_49__30_), .CO(
        u5_mult_82_CARRYB_50__29_), .S(u5_mult_82_SUMB_50__29_) );
  FA_X1 u5_mult_82_S2_50_28 ( .A(u5_mult_82_ab_50__28_), .B(
        u5_mult_82_CARRYB_49__28_), .CI(u5_mult_82_SUMB_49__29_), .CO(
        u5_mult_82_CARRYB_50__28_), .S(u5_mult_82_SUMB_50__28_) );
  FA_X1 u5_mult_82_S2_50_27 ( .A(u5_mult_82_ab_50__27_), .B(
        u5_mult_82_CARRYB_49__27_), .CI(u5_mult_82_SUMB_49__28_), .CO(
        u5_mult_82_CARRYB_50__27_), .S(u5_mult_82_SUMB_50__27_) );
  FA_X1 u5_mult_82_S2_50_26 ( .A(u5_mult_82_ab_50__26_), .B(
        u5_mult_82_CARRYB_49__26_), .CI(u5_mult_82_SUMB_49__27_), .CO(
        u5_mult_82_CARRYB_50__26_), .S(u5_mult_82_SUMB_50__26_) );
  FA_X1 u5_mult_82_S2_50_25 ( .A(u5_mult_82_ab_50__25_), .B(
        u5_mult_82_CARRYB_49__25_), .CI(u5_mult_82_SUMB_49__26_), .CO(
        u5_mult_82_CARRYB_50__25_), .S(u5_mult_82_SUMB_50__25_) );
  FA_X1 u5_mult_82_S2_50_24 ( .A(u5_mult_82_ab_50__24_), .B(
        u5_mult_82_CARRYB_49__24_), .CI(u5_mult_82_SUMB_49__25_), .CO(
        u5_mult_82_CARRYB_50__24_), .S(u5_mult_82_SUMB_50__24_) );
  FA_X1 u5_mult_82_S2_50_23 ( .A(u5_mult_82_ab_50__23_), .B(
        u5_mult_82_CARRYB_49__23_), .CI(u5_mult_82_SUMB_49__24_), .CO(
        u5_mult_82_CARRYB_50__23_), .S(u5_mult_82_SUMB_50__23_) );
  FA_X1 u5_mult_82_S2_50_22 ( .A(u5_mult_82_ab_50__22_), .B(
        u5_mult_82_CARRYB_49__22_), .CI(u5_mult_82_SUMB_49__23_), .CO(
        u5_mult_82_CARRYB_50__22_), .S(u5_mult_82_SUMB_50__22_) );
  FA_X1 u5_mult_82_S2_50_21 ( .A(u5_mult_82_ab_50__21_), .B(
        u5_mult_82_CARRYB_49__21_), .CI(u5_mult_82_SUMB_49__22_), .CO(
        u5_mult_82_CARRYB_50__21_), .S(u5_mult_82_SUMB_50__21_) );
  FA_X1 u5_mult_82_S2_50_20 ( .A(u5_mult_82_ab_50__20_), .B(
        u5_mult_82_CARRYB_49__20_), .CI(u5_mult_82_SUMB_49__21_), .CO(
        u5_mult_82_CARRYB_50__20_), .S(u5_mult_82_SUMB_50__20_) );
  FA_X1 u5_mult_82_S2_50_19 ( .A(u5_mult_82_ab_50__19_), .B(
        u5_mult_82_CARRYB_49__19_), .CI(u5_mult_82_SUMB_49__20_), .CO(
        u5_mult_82_CARRYB_50__19_), .S(u5_mult_82_SUMB_50__19_) );
  FA_X1 u5_mult_82_S2_50_18 ( .A(u5_mult_82_ab_50__18_), .B(
        u5_mult_82_CARRYB_49__18_), .CI(u5_mult_82_SUMB_49__19_), .CO(
        u5_mult_82_CARRYB_50__18_), .S(u5_mult_82_SUMB_50__18_) );
  FA_X1 u5_mult_82_S2_50_17 ( .A(u5_mult_82_ab_50__17_), .B(
        u5_mult_82_CARRYB_49__17_), .CI(u5_mult_82_SUMB_49__18_), .CO(
        u5_mult_82_CARRYB_50__17_), .S(u5_mult_82_SUMB_50__17_) );
  FA_X1 u5_mult_82_S2_50_16 ( .A(u5_mult_82_ab_50__16_), .B(
        u5_mult_82_CARRYB_49__16_), .CI(u5_mult_82_SUMB_49__17_), .CO(
        u5_mult_82_CARRYB_50__16_), .S(u5_mult_82_SUMB_50__16_) );
  FA_X1 u5_mult_82_S2_50_15 ( .A(u5_mult_82_ab_50__15_), .B(
        u5_mult_82_CARRYB_49__15_), .CI(u5_mult_82_SUMB_49__16_), .CO(
        u5_mult_82_CARRYB_50__15_), .S(u5_mult_82_SUMB_50__15_) );
  FA_X1 u5_mult_82_S2_50_14 ( .A(u5_mult_82_ab_50__14_), .B(
        u5_mult_82_CARRYB_49__14_), .CI(u5_mult_82_SUMB_49__15_), .CO(
        u5_mult_82_CARRYB_50__14_), .S(u5_mult_82_SUMB_50__14_) );
  FA_X1 u5_mult_82_S2_50_13 ( .A(u5_mult_82_ab_50__13_), .B(
        u5_mult_82_CARRYB_49__13_), .CI(u5_mult_82_SUMB_49__14_), .CO(
        u5_mult_82_CARRYB_50__13_), .S(u5_mult_82_SUMB_50__13_) );
  FA_X1 u5_mult_82_S2_50_12 ( .A(u5_mult_82_ab_50__12_), .B(
        u5_mult_82_CARRYB_49__12_), .CI(u5_mult_82_SUMB_49__13_), .CO(
        u5_mult_82_CARRYB_50__12_), .S(u5_mult_82_SUMB_50__12_) );
  FA_X1 u5_mult_82_S2_50_11 ( .A(u5_mult_82_ab_50__11_), .B(
        u5_mult_82_CARRYB_49__11_), .CI(u5_mult_82_SUMB_49__12_), .CO(
        u5_mult_82_CARRYB_50__11_), .S(u5_mult_82_SUMB_50__11_) );
  FA_X1 u5_mult_82_S2_50_10 ( .A(u5_mult_82_ab_50__10_), .B(
        u5_mult_82_CARRYB_49__10_), .CI(u5_mult_82_SUMB_49__11_), .CO(
        u5_mult_82_CARRYB_50__10_), .S(u5_mult_82_SUMB_50__10_) );
  FA_X1 u5_mult_82_S2_50_9 ( .A(u5_mult_82_ab_50__9_), .B(
        u5_mult_82_CARRYB_49__9_), .CI(u5_mult_82_SUMB_49__10_), .CO(
        u5_mult_82_CARRYB_50__9_), .S(u5_mult_82_SUMB_50__9_) );
  FA_X1 u5_mult_82_S2_50_8 ( .A(u5_mult_82_ab_50__8_), .B(
        u5_mult_82_CARRYB_49__8_), .CI(u5_mult_82_SUMB_49__9_), .CO(
        u5_mult_82_CARRYB_50__8_), .S(u5_mult_82_SUMB_50__8_) );
  FA_X1 u5_mult_82_S2_50_7 ( .A(u5_mult_82_ab_50__7_), .B(
        u5_mult_82_CARRYB_49__7_), .CI(u5_mult_82_SUMB_49__8_), .CO(
        u5_mult_82_CARRYB_50__7_), .S(u5_mult_82_SUMB_50__7_) );
  FA_X1 u5_mult_82_S2_50_6 ( .A(u5_mult_82_ab_50__6_), .B(
        u5_mult_82_CARRYB_49__6_), .CI(u5_mult_82_SUMB_49__7_), .CO(
        u5_mult_82_CARRYB_50__6_), .S(u5_mult_82_SUMB_50__6_) );
  FA_X1 u5_mult_82_S2_50_5 ( .A(u5_mult_82_ab_50__5_), .B(
        u5_mult_82_CARRYB_49__5_), .CI(u5_mult_82_SUMB_49__6_), .CO(
        u5_mult_82_CARRYB_50__5_), .S(u5_mult_82_SUMB_50__5_) );
  FA_X1 u5_mult_82_S2_50_4 ( .A(u5_mult_82_ab_50__4_), .B(
        u5_mult_82_CARRYB_49__4_), .CI(u5_mult_82_SUMB_49__5_), .CO(
        u5_mult_82_CARRYB_50__4_), .S(u5_mult_82_SUMB_50__4_) );
  FA_X1 u5_mult_82_S2_50_3 ( .A(u5_mult_82_ab_50__3_), .B(
        u5_mult_82_CARRYB_49__3_), .CI(u5_mult_82_SUMB_49__4_), .CO(
        u5_mult_82_CARRYB_50__3_), .S(u5_mult_82_SUMB_50__3_) );
  FA_X1 u5_mult_82_S2_50_2 ( .A(u5_mult_82_ab_50__2_), .B(
        u5_mult_82_CARRYB_49__2_), .CI(u5_mult_82_SUMB_49__3_), .CO(
        u5_mult_82_CARRYB_50__2_), .S(u5_mult_82_SUMB_50__2_) );
  FA_X1 u5_mult_82_S2_50_1 ( .A(u5_mult_82_ab_50__1_), .B(
        u5_mult_82_CARRYB_49__1_), .CI(u5_mult_82_SUMB_49__2_), .CO(
        u5_mult_82_CARRYB_50__1_), .S(u5_mult_82_SUMB_50__1_) );
  FA_X1 u5_mult_82_S1_50_0 ( .A(u5_mult_82_ab_50__0_), .B(
        u5_mult_82_CARRYB_49__0_), .CI(u5_mult_82_SUMB_49__1_), .CO(
        u5_mult_82_CARRYB_50__0_), .S(u5_N50) );
  FA_X1 u5_mult_82_S3_51_51 ( .A(u5_mult_82_ab_51__51_), .B(
        u5_mult_82_CARRYB_50__51_), .CI(u5_mult_82_ab_50__52_), .CO(
        u5_mult_82_CARRYB_51__51_), .S(u5_mult_82_SUMB_51__51_) );
  FA_X1 u5_mult_82_S2_51_50 ( .A(u5_mult_82_ab_51__50_), .B(
        u5_mult_82_CARRYB_50__50_), .CI(u5_mult_82_SUMB_50__51_), .CO(
        u5_mult_82_CARRYB_51__50_), .S(u5_mult_82_SUMB_51__50_) );
  FA_X1 u5_mult_82_S2_51_49 ( .A(u5_mult_82_ab_51__49_), .B(
        u5_mult_82_CARRYB_50__49_), .CI(u5_mult_82_SUMB_50__50_), .CO(
        u5_mult_82_CARRYB_51__49_), .S(u5_mult_82_SUMB_51__49_) );
  FA_X1 u5_mult_82_S2_51_48 ( .A(u5_mult_82_ab_51__48_), .B(
        u5_mult_82_CARRYB_50__48_), .CI(u5_mult_82_SUMB_50__49_), .CO(
        u5_mult_82_CARRYB_51__48_), .S(u5_mult_82_SUMB_51__48_) );
  FA_X1 u5_mult_82_S2_51_47 ( .A(u5_mult_82_ab_51__47_), .B(
        u5_mult_82_CARRYB_50__47_), .CI(u5_mult_82_SUMB_50__48_), .CO(
        u5_mult_82_CARRYB_51__47_), .S(u5_mult_82_SUMB_51__47_) );
  FA_X1 u5_mult_82_S2_51_46 ( .A(u5_mult_82_ab_51__46_), .B(
        u5_mult_82_CARRYB_50__46_), .CI(u5_mult_82_SUMB_50__47_), .CO(
        u5_mult_82_CARRYB_51__46_), .S(u5_mult_82_SUMB_51__46_) );
  FA_X1 u5_mult_82_S2_51_45 ( .A(u5_mult_82_ab_51__45_), .B(
        u5_mult_82_CARRYB_50__45_), .CI(u5_mult_82_SUMB_50__46_), .CO(
        u5_mult_82_CARRYB_51__45_), .S(u5_mult_82_SUMB_51__45_) );
  FA_X1 u5_mult_82_S2_51_44 ( .A(u5_mult_82_ab_51__44_), .B(
        u5_mult_82_CARRYB_50__44_), .CI(u5_mult_82_SUMB_50__45_), .CO(
        u5_mult_82_CARRYB_51__44_), .S(u5_mult_82_SUMB_51__44_) );
  FA_X1 u5_mult_82_S2_51_43 ( .A(u5_mult_82_ab_51__43_), .B(
        u5_mult_82_CARRYB_50__43_), .CI(u5_mult_82_SUMB_50__44_), .CO(
        u5_mult_82_CARRYB_51__43_), .S(u5_mult_82_SUMB_51__43_) );
  FA_X1 u5_mult_82_S2_51_42 ( .A(u5_mult_82_ab_51__42_), .B(
        u5_mult_82_CARRYB_50__42_), .CI(u5_mult_82_SUMB_50__43_), .CO(
        u5_mult_82_CARRYB_51__42_), .S(u5_mult_82_SUMB_51__42_) );
  FA_X1 u5_mult_82_S2_51_41 ( .A(u5_mult_82_ab_51__41_), .B(
        u5_mult_82_CARRYB_50__41_), .CI(u5_mult_82_SUMB_50__42_), .CO(
        u5_mult_82_CARRYB_51__41_), .S(u5_mult_82_SUMB_51__41_) );
  FA_X1 u5_mult_82_S2_51_40 ( .A(u5_mult_82_ab_51__40_), .B(
        u5_mult_82_CARRYB_50__40_), .CI(u5_mult_82_SUMB_50__41_), .CO(
        u5_mult_82_CARRYB_51__40_), .S(u5_mult_82_SUMB_51__40_) );
  FA_X1 u5_mult_82_S2_51_39 ( .A(u5_mult_82_ab_51__39_), .B(
        u5_mult_82_CARRYB_50__39_), .CI(u5_mult_82_SUMB_50__40_), .CO(
        u5_mult_82_CARRYB_51__39_), .S(u5_mult_82_SUMB_51__39_) );
  FA_X1 u5_mult_82_S2_51_38 ( .A(u5_mult_82_ab_51__38_), .B(
        u5_mult_82_CARRYB_50__38_), .CI(u5_mult_82_SUMB_50__39_), .CO(
        u5_mult_82_CARRYB_51__38_), .S(u5_mult_82_SUMB_51__38_) );
  FA_X1 u5_mult_82_S2_51_37 ( .A(u5_mult_82_ab_51__37_), .B(
        u5_mult_82_CARRYB_50__37_), .CI(u5_mult_82_SUMB_50__38_), .CO(
        u5_mult_82_CARRYB_51__37_), .S(u5_mult_82_SUMB_51__37_) );
  FA_X1 u5_mult_82_S2_51_36 ( .A(u5_mult_82_ab_51__36_), .B(
        u5_mult_82_CARRYB_50__36_), .CI(u5_mult_82_SUMB_50__37_), .CO(
        u5_mult_82_CARRYB_51__36_), .S(u5_mult_82_SUMB_51__36_) );
  FA_X1 u5_mult_82_S2_51_35 ( .A(u5_mult_82_ab_51__35_), .B(
        u5_mult_82_CARRYB_50__35_), .CI(u5_mult_82_SUMB_50__36_), .CO(
        u5_mult_82_CARRYB_51__35_), .S(u5_mult_82_SUMB_51__35_) );
  FA_X1 u5_mult_82_S2_51_34 ( .A(u5_mult_82_ab_51__34_), .B(
        u5_mult_82_CARRYB_50__34_), .CI(u5_mult_82_SUMB_50__35_), .CO(
        u5_mult_82_CARRYB_51__34_), .S(u5_mult_82_SUMB_51__34_) );
  FA_X1 u5_mult_82_S2_51_33 ( .A(u5_mult_82_ab_51__33_), .B(
        u5_mult_82_CARRYB_50__33_), .CI(u5_mult_82_SUMB_50__34_), .CO(
        u5_mult_82_CARRYB_51__33_), .S(u5_mult_82_SUMB_51__33_) );
  FA_X1 u5_mult_82_S2_51_32 ( .A(u5_mult_82_ab_51__32_), .B(
        u5_mult_82_CARRYB_50__32_), .CI(u5_mult_82_SUMB_50__33_), .CO(
        u5_mult_82_CARRYB_51__32_), .S(u5_mult_82_SUMB_51__32_) );
  FA_X1 u5_mult_82_S2_51_31 ( .A(u5_mult_82_ab_51__31_), .B(
        u5_mult_82_CARRYB_50__31_), .CI(u5_mult_82_SUMB_50__32_), .CO(
        u5_mult_82_CARRYB_51__31_), .S(u5_mult_82_SUMB_51__31_) );
  FA_X1 u5_mult_82_S2_51_30 ( .A(u5_mult_82_ab_51__30_), .B(
        u5_mult_82_CARRYB_50__30_), .CI(u5_mult_82_SUMB_50__31_), .CO(
        u5_mult_82_CARRYB_51__30_), .S(u5_mult_82_SUMB_51__30_) );
  FA_X1 u5_mult_82_S2_51_29 ( .A(u5_mult_82_ab_51__29_), .B(
        u5_mult_82_CARRYB_50__29_), .CI(u5_mult_82_SUMB_50__30_), .CO(
        u5_mult_82_CARRYB_51__29_), .S(u5_mult_82_SUMB_51__29_) );
  FA_X1 u5_mult_82_S2_51_28 ( .A(u5_mult_82_ab_51__28_), .B(
        u5_mult_82_CARRYB_50__28_), .CI(u5_mult_82_SUMB_50__29_), .CO(
        u5_mult_82_CARRYB_51__28_), .S(u5_mult_82_SUMB_51__28_) );
  FA_X1 u5_mult_82_S2_51_27 ( .A(u5_mult_82_ab_51__27_), .B(
        u5_mult_82_CARRYB_50__27_), .CI(u5_mult_82_SUMB_50__28_), .CO(
        u5_mult_82_CARRYB_51__27_), .S(u5_mult_82_SUMB_51__27_) );
  FA_X1 u5_mult_82_S2_51_26 ( .A(u5_mult_82_ab_51__26_), .B(
        u5_mult_82_CARRYB_50__26_), .CI(u5_mult_82_SUMB_50__27_), .CO(
        u5_mult_82_CARRYB_51__26_), .S(u5_mult_82_SUMB_51__26_) );
  FA_X1 u5_mult_82_S2_51_25 ( .A(u5_mult_82_ab_51__25_), .B(
        u5_mult_82_CARRYB_50__25_), .CI(u5_mult_82_SUMB_50__26_), .CO(
        u5_mult_82_CARRYB_51__25_), .S(u5_mult_82_SUMB_51__25_) );
  FA_X1 u5_mult_82_S2_51_24 ( .A(u5_mult_82_ab_51__24_), .B(
        u5_mult_82_CARRYB_50__24_), .CI(u5_mult_82_SUMB_50__25_), .CO(
        u5_mult_82_CARRYB_51__24_), .S(u5_mult_82_SUMB_51__24_) );
  FA_X1 u5_mult_82_S2_51_23 ( .A(u5_mult_82_ab_51__23_), .B(
        u5_mult_82_CARRYB_50__23_), .CI(u5_mult_82_SUMB_50__24_), .CO(
        u5_mult_82_CARRYB_51__23_), .S(u5_mult_82_SUMB_51__23_) );
  FA_X1 u5_mult_82_S2_51_22 ( .A(u5_mult_82_ab_51__22_), .B(
        u5_mult_82_CARRYB_50__22_), .CI(u5_mult_82_SUMB_50__23_), .CO(
        u5_mult_82_CARRYB_51__22_), .S(u5_mult_82_SUMB_51__22_) );
  FA_X1 u5_mult_82_S2_51_21 ( .A(u5_mult_82_ab_51__21_), .B(
        u5_mult_82_CARRYB_50__21_), .CI(u5_mult_82_SUMB_50__22_), .CO(
        u5_mult_82_CARRYB_51__21_), .S(u5_mult_82_SUMB_51__21_) );
  FA_X1 u5_mult_82_S2_51_20 ( .A(u5_mult_82_ab_51__20_), .B(
        u5_mult_82_CARRYB_50__20_), .CI(u5_mult_82_SUMB_50__21_), .CO(
        u5_mult_82_CARRYB_51__20_), .S(u5_mult_82_SUMB_51__20_) );
  FA_X1 u5_mult_82_S2_51_19 ( .A(u5_mult_82_ab_51__19_), .B(
        u5_mult_82_CARRYB_50__19_), .CI(u5_mult_82_SUMB_50__20_), .CO(
        u5_mult_82_CARRYB_51__19_), .S(u5_mult_82_SUMB_51__19_) );
  FA_X1 u5_mult_82_S2_51_18 ( .A(u5_mult_82_ab_51__18_), .B(
        u5_mult_82_CARRYB_50__18_), .CI(u5_mult_82_SUMB_50__19_), .CO(
        u5_mult_82_CARRYB_51__18_), .S(u5_mult_82_SUMB_51__18_) );
  FA_X1 u5_mult_82_S2_51_17 ( .A(u5_mult_82_ab_51__17_), .B(
        u5_mult_82_CARRYB_50__17_), .CI(u5_mult_82_SUMB_50__18_), .CO(
        u5_mult_82_CARRYB_51__17_), .S(u5_mult_82_SUMB_51__17_) );
  FA_X1 u5_mult_82_S2_51_16 ( .A(u5_mult_82_ab_51__16_), .B(
        u5_mult_82_CARRYB_50__16_), .CI(u5_mult_82_SUMB_50__17_), .CO(
        u5_mult_82_CARRYB_51__16_), .S(u5_mult_82_SUMB_51__16_) );
  FA_X1 u5_mult_82_S2_51_15 ( .A(u5_mult_82_ab_51__15_), .B(
        u5_mult_82_CARRYB_50__15_), .CI(u5_mult_82_SUMB_50__16_), .CO(
        u5_mult_82_CARRYB_51__15_), .S(u5_mult_82_SUMB_51__15_) );
  FA_X1 u5_mult_82_S2_51_14 ( .A(u5_mult_82_ab_51__14_), .B(
        u5_mult_82_CARRYB_50__14_), .CI(u5_mult_82_SUMB_50__15_), .CO(
        u5_mult_82_CARRYB_51__14_), .S(u5_mult_82_SUMB_51__14_) );
  FA_X1 u5_mult_82_S2_51_13 ( .A(u5_mult_82_ab_51__13_), .B(
        u5_mult_82_CARRYB_50__13_), .CI(u5_mult_82_SUMB_50__14_), .CO(
        u5_mult_82_CARRYB_51__13_), .S(u5_mult_82_SUMB_51__13_) );
  FA_X1 u5_mult_82_S2_51_12 ( .A(u5_mult_82_ab_51__12_), .B(
        u5_mult_82_CARRYB_50__12_), .CI(u5_mult_82_SUMB_50__13_), .CO(
        u5_mult_82_CARRYB_51__12_), .S(u5_mult_82_SUMB_51__12_) );
  FA_X1 u5_mult_82_S2_51_11 ( .A(u5_mult_82_ab_51__11_), .B(
        u5_mult_82_CARRYB_50__11_), .CI(u5_mult_82_SUMB_50__12_), .CO(
        u5_mult_82_CARRYB_51__11_), .S(u5_mult_82_SUMB_51__11_) );
  FA_X1 u5_mult_82_S2_51_10 ( .A(u5_mult_82_ab_51__10_), .B(
        u5_mult_82_CARRYB_50__10_), .CI(u5_mult_82_SUMB_50__11_), .CO(
        u5_mult_82_CARRYB_51__10_), .S(u5_mult_82_SUMB_51__10_) );
  FA_X1 u5_mult_82_S2_51_9 ( .A(u5_mult_82_ab_51__9_), .B(
        u5_mult_82_CARRYB_50__9_), .CI(u5_mult_82_SUMB_50__10_), .CO(
        u5_mult_82_CARRYB_51__9_), .S(u5_mult_82_SUMB_51__9_) );
  FA_X1 u5_mult_82_S2_51_8 ( .A(u5_mult_82_ab_51__8_), .B(
        u5_mult_82_CARRYB_50__8_), .CI(u5_mult_82_SUMB_50__9_), .CO(
        u5_mult_82_CARRYB_51__8_), .S(u5_mult_82_SUMB_51__8_) );
  FA_X1 u5_mult_82_S2_51_7 ( .A(u5_mult_82_ab_51__7_), .B(
        u5_mult_82_CARRYB_50__7_), .CI(u5_mult_82_SUMB_50__8_), .CO(
        u5_mult_82_CARRYB_51__7_), .S(u5_mult_82_SUMB_51__7_) );
  FA_X1 u5_mult_82_S2_51_6 ( .A(u5_mult_82_ab_51__6_), .B(
        u5_mult_82_CARRYB_50__6_), .CI(u5_mult_82_SUMB_50__7_), .CO(
        u5_mult_82_CARRYB_51__6_), .S(u5_mult_82_SUMB_51__6_) );
  FA_X1 u5_mult_82_S2_51_5 ( .A(u5_mult_82_ab_51__5_), .B(
        u5_mult_82_CARRYB_50__5_), .CI(u5_mult_82_SUMB_50__6_), .CO(
        u5_mult_82_CARRYB_51__5_), .S(u5_mult_82_SUMB_51__5_) );
  FA_X1 u5_mult_82_S2_51_4 ( .A(u5_mult_82_ab_51__4_), .B(
        u5_mult_82_CARRYB_50__4_), .CI(u5_mult_82_SUMB_50__5_), .CO(
        u5_mult_82_CARRYB_51__4_), .S(u5_mult_82_SUMB_51__4_) );
  FA_X1 u5_mult_82_S2_51_3 ( .A(u5_mult_82_ab_51__3_), .B(
        u5_mult_82_CARRYB_50__3_), .CI(u5_mult_82_SUMB_50__4_), .CO(
        u5_mult_82_CARRYB_51__3_), .S(u5_mult_82_SUMB_51__3_) );
  FA_X1 u5_mult_82_S2_51_2 ( .A(u5_mult_82_ab_51__2_), .B(
        u5_mult_82_CARRYB_50__2_), .CI(u5_mult_82_SUMB_50__3_), .CO(
        u5_mult_82_CARRYB_51__2_), .S(u5_mult_82_SUMB_51__2_) );
  FA_X1 u5_mult_82_S2_51_1 ( .A(u5_mult_82_ab_51__1_), .B(
        u5_mult_82_CARRYB_50__1_), .CI(u5_mult_82_SUMB_50__2_), .CO(
        u5_mult_82_CARRYB_51__1_), .S(u5_mult_82_SUMB_51__1_) );
  FA_X1 u5_mult_82_S1_51_0 ( .A(u5_mult_82_ab_51__0_), .B(
        u5_mult_82_CARRYB_50__0_), .CI(u5_mult_82_SUMB_50__1_), .CO(
        u5_mult_82_CARRYB_51__0_), .S(u5_N51) );
  FA_X1 u5_mult_82_S5_51 ( .A(u5_mult_82_ab_52__51_), .B(
        u5_mult_82_CARRYB_51__51_), .CI(u5_mult_82_ab_51__52_), .CO(
        u5_mult_82_CARRYB_52__51_), .S(u5_mult_82_SUMB_52__51_) );
  FA_X1 u5_mult_82_S4_50 ( .A(u5_mult_82_ab_52__50_), .B(
        u5_mult_82_CARRYB_51__50_), .CI(u5_mult_82_SUMB_51__51_), .CO(
        u5_mult_82_CARRYB_52__50_), .S(u5_mult_82_SUMB_52__50_) );
  FA_X1 u5_mult_82_S4_49 ( .A(u5_mult_82_ab_52__49_), .B(
        u5_mult_82_CARRYB_51__49_), .CI(u5_mult_82_SUMB_51__50_), .CO(
        u5_mult_82_CARRYB_52__49_), .S(u5_mult_82_SUMB_52__49_) );
  FA_X1 u5_mult_82_S4_48 ( .A(u5_mult_82_ab_52__48_), .B(
        u5_mult_82_CARRYB_51__48_), .CI(u5_mult_82_SUMB_51__49_), .CO(
        u5_mult_82_CARRYB_52__48_), .S(u5_mult_82_SUMB_52__48_) );
  FA_X1 u5_mult_82_S4_47 ( .A(u5_mult_82_ab_52__47_), .B(
        u5_mult_82_CARRYB_51__47_), .CI(u5_mult_82_SUMB_51__48_), .CO(
        u5_mult_82_CARRYB_52__47_), .S(u5_mult_82_SUMB_52__47_) );
  FA_X1 u5_mult_82_S4_46 ( .A(u5_mult_82_ab_52__46_), .B(
        u5_mult_82_CARRYB_51__46_), .CI(u5_mult_82_SUMB_51__47_), .CO(
        u5_mult_82_CARRYB_52__46_), .S(u5_mult_82_SUMB_52__46_) );
  FA_X1 u5_mult_82_S4_45 ( .A(u5_mult_82_ab_52__45_), .B(
        u5_mult_82_CARRYB_51__45_), .CI(u5_mult_82_SUMB_51__46_), .CO(
        u5_mult_82_CARRYB_52__45_), .S(u5_mult_82_SUMB_52__45_) );
  FA_X1 u5_mult_82_S4_44 ( .A(u5_mult_82_ab_52__44_), .B(
        u5_mult_82_CARRYB_51__44_), .CI(u5_mult_82_SUMB_51__45_), .CO(
        u5_mult_82_CARRYB_52__44_), .S(u5_mult_82_SUMB_52__44_) );
  FA_X1 u5_mult_82_S4_43 ( .A(u5_mult_82_ab_52__43_), .B(
        u5_mult_82_CARRYB_51__43_), .CI(u5_mult_82_SUMB_51__44_), .CO(
        u5_mult_82_CARRYB_52__43_), .S(u5_mult_82_SUMB_52__43_) );
  FA_X1 u5_mult_82_S4_42 ( .A(u5_mult_82_ab_52__42_), .B(
        u5_mult_82_CARRYB_51__42_), .CI(u5_mult_82_SUMB_51__43_), .CO(
        u5_mult_82_CARRYB_52__42_), .S(u5_mult_82_SUMB_52__42_) );
  FA_X1 u5_mult_82_S4_41 ( .A(u5_mult_82_ab_52__41_), .B(
        u5_mult_82_CARRYB_51__41_), .CI(u5_mult_82_SUMB_51__42_), .CO(
        u5_mult_82_CARRYB_52__41_), .S(u5_mult_82_SUMB_52__41_) );
  FA_X1 u5_mult_82_S4_40 ( .A(u5_mult_82_ab_52__40_), .B(
        u5_mult_82_CARRYB_51__40_), .CI(u5_mult_82_SUMB_51__41_), .CO(
        u5_mult_82_CARRYB_52__40_), .S(u5_mult_82_SUMB_52__40_) );
  FA_X1 u5_mult_82_S4_39 ( .A(u5_mult_82_ab_52__39_), .B(
        u5_mult_82_CARRYB_51__39_), .CI(u5_mult_82_SUMB_51__40_), .CO(
        u5_mult_82_CARRYB_52__39_), .S(u5_mult_82_SUMB_52__39_) );
  FA_X1 u5_mult_82_S4_38 ( .A(u5_mult_82_ab_52__38_), .B(
        u5_mult_82_CARRYB_51__38_), .CI(u5_mult_82_SUMB_51__39_), .CO(
        u5_mult_82_CARRYB_52__38_), .S(u5_mult_82_SUMB_52__38_) );
  FA_X1 u5_mult_82_S4_37 ( .A(u5_mult_82_ab_52__37_), .B(
        u5_mult_82_CARRYB_51__37_), .CI(u5_mult_82_SUMB_51__38_), .CO(
        u5_mult_82_CARRYB_52__37_), .S(u5_mult_82_SUMB_52__37_) );
  FA_X1 u5_mult_82_S4_36 ( .A(u5_mult_82_ab_52__36_), .B(
        u5_mult_82_CARRYB_51__36_), .CI(u5_mult_82_SUMB_51__37_), .CO(
        u5_mult_82_CARRYB_52__36_), .S(u5_mult_82_SUMB_52__36_) );
  FA_X1 u5_mult_82_S4_35 ( .A(u5_mult_82_ab_52__35_), .B(
        u5_mult_82_CARRYB_51__35_), .CI(u5_mult_82_SUMB_51__36_), .CO(
        u5_mult_82_CARRYB_52__35_), .S(u5_mult_82_SUMB_52__35_) );
  FA_X1 u5_mult_82_S4_34 ( .A(u5_mult_82_ab_52__34_), .B(
        u5_mult_82_CARRYB_51__34_), .CI(u5_mult_82_SUMB_51__35_), .CO(
        u5_mult_82_CARRYB_52__34_), .S(u5_mult_82_SUMB_52__34_) );
  FA_X1 u5_mult_82_S4_33 ( .A(u5_mult_82_ab_52__33_), .B(
        u5_mult_82_CARRYB_51__33_), .CI(u5_mult_82_SUMB_51__34_), .CO(
        u5_mult_82_CARRYB_52__33_), .S(u5_mult_82_SUMB_52__33_) );
  FA_X1 u5_mult_82_S4_32 ( .A(u5_mult_82_ab_52__32_), .B(
        u5_mult_82_CARRYB_51__32_), .CI(u5_mult_82_SUMB_51__33_), .CO(
        u5_mult_82_CARRYB_52__32_), .S(u5_mult_82_SUMB_52__32_) );
  FA_X1 u5_mult_82_S4_31 ( .A(u5_mult_82_ab_52__31_), .B(
        u5_mult_82_CARRYB_51__31_), .CI(u5_mult_82_SUMB_51__32_), .CO(
        u5_mult_82_CARRYB_52__31_), .S(u5_mult_82_SUMB_52__31_) );
  FA_X1 u5_mult_82_S4_30 ( .A(u5_mult_82_ab_52__30_), .B(
        u5_mult_82_CARRYB_51__30_), .CI(u5_mult_82_SUMB_51__31_), .CO(
        u5_mult_82_CARRYB_52__30_), .S(u5_mult_82_SUMB_52__30_) );
  FA_X1 u5_mult_82_S4_29 ( .A(u5_mult_82_ab_52__29_), .B(
        u5_mult_82_CARRYB_51__29_), .CI(u5_mult_82_SUMB_51__30_), .CO(
        u5_mult_82_CARRYB_52__29_), .S(u5_mult_82_SUMB_52__29_) );
  FA_X1 u5_mult_82_S4_28 ( .A(u5_mult_82_ab_52__28_), .B(
        u5_mult_82_CARRYB_51__28_), .CI(u5_mult_82_SUMB_51__29_), .CO(
        u5_mult_82_CARRYB_52__28_), .S(u5_mult_82_SUMB_52__28_) );
  FA_X1 u5_mult_82_S4_27 ( .A(u5_mult_82_ab_52__27_), .B(
        u5_mult_82_CARRYB_51__27_), .CI(u5_mult_82_SUMB_51__28_), .CO(
        u5_mult_82_CARRYB_52__27_), .S(u5_mult_82_SUMB_52__27_) );
  FA_X1 u5_mult_82_S4_26 ( .A(u5_mult_82_ab_52__26_), .B(
        u5_mult_82_CARRYB_51__26_), .CI(u5_mult_82_SUMB_51__27_), .CO(
        u5_mult_82_CARRYB_52__26_), .S(u5_mult_82_SUMB_52__26_) );
  FA_X1 u5_mult_82_S4_25 ( .A(u5_mult_82_ab_52__25_), .B(
        u5_mult_82_CARRYB_51__25_), .CI(u5_mult_82_SUMB_51__26_), .CO(
        u5_mult_82_CARRYB_52__25_), .S(u5_mult_82_SUMB_52__25_) );
  FA_X1 u5_mult_82_S4_24 ( .A(u5_mult_82_ab_52__24_), .B(
        u5_mult_82_CARRYB_51__24_), .CI(u5_mult_82_SUMB_51__25_), .CO(
        u5_mult_82_CARRYB_52__24_), .S(u5_mult_82_SUMB_52__24_) );
  FA_X1 u5_mult_82_S4_23 ( .A(u5_mult_82_ab_52__23_), .B(
        u5_mult_82_CARRYB_51__23_), .CI(u5_mult_82_SUMB_51__24_), .CO(
        u5_mult_82_CARRYB_52__23_), .S(u5_mult_82_SUMB_52__23_) );
  FA_X1 u5_mult_82_S4_22 ( .A(u5_mult_82_ab_52__22_), .B(
        u5_mult_82_CARRYB_51__22_), .CI(u5_mult_82_SUMB_51__23_), .CO(
        u5_mult_82_CARRYB_52__22_), .S(u5_mult_82_SUMB_52__22_) );
  FA_X1 u5_mult_82_S4_21 ( .A(u5_mult_82_ab_52__21_), .B(
        u5_mult_82_CARRYB_51__21_), .CI(u5_mult_82_SUMB_51__22_), .CO(
        u5_mult_82_CARRYB_52__21_), .S(u5_mult_82_SUMB_52__21_) );
  FA_X1 u5_mult_82_S4_20 ( .A(u5_mult_82_ab_52__20_), .B(
        u5_mult_82_CARRYB_51__20_), .CI(u5_mult_82_SUMB_51__21_), .CO(
        u5_mult_82_CARRYB_52__20_), .S(u5_mult_82_SUMB_52__20_) );
  FA_X1 u5_mult_82_S4_19 ( .A(u5_mult_82_ab_52__19_), .B(
        u5_mult_82_CARRYB_51__19_), .CI(u5_mult_82_SUMB_51__20_), .CO(
        u5_mult_82_CARRYB_52__19_), .S(u5_mult_82_SUMB_52__19_) );
  FA_X1 u5_mult_82_S4_18 ( .A(u5_mult_82_ab_52__18_), .B(
        u5_mult_82_CARRYB_51__18_), .CI(u5_mult_82_SUMB_51__19_), .CO(
        u5_mult_82_CARRYB_52__18_), .S(u5_mult_82_SUMB_52__18_) );
  FA_X1 u5_mult_82_S4_17 ( .A(u5_mult_82_ab_52__17_), .B(
        u5_mult_82_CARRYB_51__17_), .CI(u5_mult_82_SUMB_51__18_), .CO(
        u5_mult_82_CARRYB_52__17_), .S(u5_mult_82_SUMB_52__17_) );
  FA_X1 u5_mult_82_S4_16 ( .A(u5_mult_82_ab_52__16_), .B(
        u5_mult_82_CARRYB_51__16_), .CI(u5_mult_82_SUMB_51__17_), .CO(
        u5_mult_82_CARRYB_52__16_), .S(u5_mult_82_SUMB_52__16_) );
  FA_X1 u5_mult_82_S4_15 ( .A(u5_mult_82_ab_52__15_), .B(
        u5_mult_82_CARRYB_51__15_), .CI(u5_mult_82_SUMB_51__16_), .CO(
        u5_mult_82_CARRYB_52__15_), .S(u5_mult_82_SUMB_52__15_) );
  FA_X1 u5_mult_82_S4_14 ( .A(u5_mult_82_ab_52__14_), .B(
        u5_mult_82_CARRYB_51__14_), .CI(u5_mult_82_SUMB_51__15_), .CO(
        u5_mult_82_CARRYB_52__14_), .S(u5_mult_82_SUMB_52__14_) );
  FA_X1 u5_mult_82_S4_13 ( .A(u5_mult_82_ab_52__13_), .B(
        u5_mult_82_CARRYB_51__13_), .CI(u5_mult_82_SUMB_51__14_), .CO(
        u5_mult_82_CARRYB_52__13_), .S(u5_mult_82_SUMB_52__13_) );
  FA_X1 u5_mult_82_S4_12 ( .A(u5_mult_82_ab_52__12_), .B(
        u5_mult_82_CARRYB_51__12_), .CI(u5_mult_82_SUMB_51__13_), .CO(
        u5_mult_82_CARRYB_52__12_), .S(u5_mult_82_SUMB_52__12_) );
  FA_X1 u5_mult_82_S4_11 ( .A(u5_mult_82_ab_52__11_), .B(
        u5_mult_82_CARRYB_51__11_), .CI(u5_mult_82_SUMB_51__12_), .CO(
        u5_mult_82_CARRYB_52__11_), .S(u5_mult_82_SUMB_52__11_) );
  FA_X1 u5_mult_82_S4_10 ( .A(u5_mult_82_ab_52__10_), .B(
        u5_mult_82_CARRYB_51__10_), .CI(u5_mult_82_SUMB_51__11_), .CO(
        u5_mult_82_CARRYB_52__10_), .S(u5_mult_82_SUMB_52__10_) );
  FA_X1 u5_mult_82_S4_9 ( .A(u5_mult_82_ab_52__9_), .B(
        u5_mult_82_CARRYB_51__9_), .CI(u5_mult_82_SUMB_51__10_), .CO(
        u5_mult_82_CARRYB_52__9_), .S(u5_mult_82_SUMB_52__9_) );
  FA_X1 u5_mult_82_S4_8 ( .A(u5_mult_82_ab_52__8_), .B(
        u5_mult_82_CARRYB_51__8_), .CI(u5_mult_82_SUMB_51__9_), .CO(
        u5_mult_82_CARRYB_52__8_), .S(u5_mult_82_SUMB_52__8_) );
  FA_X1 u5_mult_82_S4_7 ( .A(u5_mult_82_ab_52__7_), .B(
        u5_mult_82_CARRYB_51__7_), .CI(u5_mult_82_SUMB_51__8_), .CO(
        u5_mult_82_CARRYB_52__7_), .S(u5_mult_82_SUMB_52__7_) );
  FA_X1 u5_mult_82_S4_6 ( .A(u5_mult_82_ab_52__6_), .B(
        u5_mult_82_CARRYB_51__6_), .CI(u5_mult_82_SUMB_51__7_), .CO(
        u5_mult_82_CARRYB_52__6_), .S(u5_mult_82_SUMB_52__6_) );
  FA_X1 u5_mult_82_S4_5 ( .A(u5_mult_82_ab_52__5_), .B(
        u5_mult_82_CARRYB_51__5_), .CI(u5_mult_82_SUMB_51__6_), .CO(
        u5_mult_82_CARRYB_52__5_), .S(u5_mult_82_SUMB_52__5_) );
  FA_X1 u5_mult_82_S4_4 ( .A(u5_mult_82_ab_52__4_), .B(
        u5_mult_82_CARRYB_51__4_), .CI(u5_mult_82_SUMB_51__5_), .CO(
        u5_mult_82_CARRYB_52__4_), .S(u5_mult_82_SUMB_52__4_) );
  FA_X1 u5_mult_82_S4_3 ( .A(u5_mult_82_ab_52__3_), .B(
        u5_mult_82_CARRYB_51__3_), .CI(u5_mult_82_SUMB_51__4_), .CO(
        u5_mult_82_CARRYB_52__3_), .S(u5_mult_82_SUMB_52__3_) );
  FA_X1 u5_mult_82_S4_2 ( .A(u5_mult_82_ab_52__2_), .B(
        u5_mult_82_CARRYB_51__2_), .CI(u5_mult_82_SUMB_51__3_), .CO(
        u5_mult_82_CARRYB_52__2_), .S(u5_mult_82_SUMB_52__2_) );
  FA_X1 u5_mult_82_S4_1 ( .A(u5_mult_82_ab_52__1_), .B(
        u5_mult_82_CARRYB_51__1_), .CI(u5_mult_82_SUMB_51__2_), .CO(
        u5_mult_82_CARRYB_52__1_), .S(u5_mult_82_SUMB_52__1_) );
  FA_X1 u5_mult_82_S4_0 ( .A(u5_mult_82_ab_52__0_), .B(
        u5_mult_82_CARRYB_51__0_), .CI(u5_mult_82_SUMB_51__1_), .CO(
        u5_mult_82_CARRYB_52__0_), .S(u5_N52) );
  NOR2_X1 u5_mult_82_FS_1_U357 ( .A1(u5_mult_82_n206), .A2(u5_mult_82_n104), 
        .ZN(u5_mult_82_FS_1_n274) );
  NAND2_X1 u5_mult_82_FS_1_U356 ( .A1(u5_mult_82_n206), .A2(u5_mult_82_n104), 
        .ZN(u5_mult_82_FS_1_n276) );
  NAND2_X1 u5_mult_82_FS_1_U355 ( .A1(u5_mult_82_FS_1_n5), .A2(
        u5_mult_82_FS_1_n276), .ZN(u5_mult_82_FS_1_n277) );
  NOR2_X1 u5_mult_82_FS_1_U354 ( .A1(u5_mult_82_n205), .A2(u5_mult_82_n103), 
        .ZN(u5_mult_82_FS_1_n76) );
  NOR2_X1 u5_mult_82_FS_1_U353 ( .A1(u5_mult_82_n200), .A2(u5_mult_82_n99), 
        .ZN(u5_mult_82_FS_1_n80) );
  NOR2_X1 u5_mult_82_FS_1_U352 ( .A1(u5_mult_82_n204), .A2(u5_mult_82_n102), 
        .ZN(u5_mult_82_FS_1_n90) );
  NOR2_X1 u5_mult_82_FS_1_U351 ( .A1(u5_mult_82_n203), .A2(u5_mult_82_n101), 
        .ZN(u5_mult_82_FS_1_n93) );
  NOR2_X1 u5_mult_82_FS_1_U350 ( .A1(u5_mult_82_n195), .A2(u5_mult_82_n93), 
        .ZN(u5_mult_82_FS_1_n126) );
  NOR2_X1 u5_mult_82_FS_1_U349 ( .A1(u5_mult_82_n177), .A2(u5_mult_82_n76), 
        .ZN(u5_mult_82_FS_1_n128) );
  NOR2_X1 u5_mult_82_FS_1_U348 ( .A1(u5_mult_82_n194), .A2(u5_mult_82_n92), 
        .ZN(u5_mult_82_FS_1_n129) );
  NOR2_X1 u5_mult_82_FS_1_U347 ( .A1(u5_mult_82_n193), .A2(u5_mult_82_n91), 
        .ZN(u5_mult_82_FS_1_n133) );
  NOR4_X1 u5_mult_82_FS_1_U346 ( .A1(u5_mult_82_FS_1_n126), .A2(
        u5_mult_82_FS_1_n128), .A3(u5_mult_82_FS_1_n129), .A4(
        u5_mult_82_FS_1_n133), .ZN(u5_mult_82_FS_1_n119) );
  NOR2_X1 u5_mult_82_FS_1_U345 ( .A1(u5_mult_82_n192), .A2(u5_mult_82_n90), 
        .ZN(u5_mult_82_FS_1_n289) );
  NOR2_X1 u5_mult_82_FS_1_U344 ( .A1(u5_mult_82_n191), .A2(u5_mult_82_n89), 
        .ZN(u5_mult_82_FS_1_n144) );
  NAND2_X1 u5_mult_82_FS_1_U343 ( .A1(u5_mult_82_n190), .A2(u5_mult_82_n88), 
        .ZN(u5_mult_82_FS_1_n151) );
  NAND2_X1 u5_mult_82_FS_1_U342 ( .A1(u5_mult_82_n191), .A2(u5_mult_82_n89), 
        .ZN(u5_mult_82_FS_1_n145) );
  OAI21_X1 u5_mult_82_FS_1_U341 ( .B1(u5_mult_82_FS_1_n144), .B2(
        u5_mult_82_FS_1_n151), .A(u5_mult_82_FS_1_n145), .ZN(
        u5_mult_82_FS_1_n305) );
  OR2_X1 u5_mult_82_FS_1_U340 ( .A1(u5_mult_82_n173), .A2(u5_mult_82_n77), 
        .ZN(u5_mult_82_FS_1_n141) );
  NAND2_X1 u5_mult_82_FS_1_U339 ( .A1(u5_mult_82_n173), .A2(u5_mult_82_n77), 
        .ZN(u5_mult_82_FS_1_n146) );
  AOI21_X1 u5_mult_82_FS_1_U338 ( .B1(u5_mult_82_FS_1_n305), .B2(
        u5_mult_82_FS_1_n141), .A(u5_mult_82_FS_1_n28), .ZN(
        u5_mult_82_FS_1_n304) );
  NAND2_X1 u5_mult_82_FS_1_U337 ( .A1(u5_mult_82_n192), .A2(u5_mult_82_n90), 
        .ZN(u5_mult_82_FS_1_n142) );
  OAI21_X1 u5_mult_82_FS_1_U336 ( .B1(u5_mult_82_FS_1_n289), .B2(
        u5_mult_82_FS_1_n304), .A(u5_mult_82_FS_1_n142), .ZN(
        u5_mult_82_FS_1_n136) );
  NOR2_X1 u5_mult_82_FS_1_U335 ( .A1(u5_mult_82_n190), .A2(u5_mult_82_n88), 
        .ZN(u5_mult_82_FS_1_n150) );
  NOR2_X1 u5_mult_82_FS_1_U334 ( .A1(u5_mult_82_n176), .A2(u5_mult_82_n75), 
        .ZN(u5_mult_82_FS_1_n156) );
  NOR2_X1 u5_mult_82_FS_1_U333 ( .A1(u5_mult_82_n175), .A2(u5_mult_82_n74), 
        .ZN(u5_mult_82_FS_1_n164) );
  NOR2_X1 u5_mult_82_FS_1_U332 ( .A1(u5_mult_82_n189), .A2(u5_mult_82_n87), 
        .ZN(u5_mult_82_FS_1_n298) );
  OR2_X1 u5_mult_82_FS_1_U331 ( .A1(u5_mult_82_n172), .A2(u5_mult_82_n60), 
        .ZN(u5_mult_82_FS_1_n192) );
  NOR2_X1 u5_mult_82_FS_1_U330 ( .A1(u5_mult_82_n188), .A2(u5_mult_82_n71), 
        .ZN(u5_mult_82_FS_1_n195) );
  NOR2_X1 u5_mult_82_FS_1_U329 ( .A1(u5_mult_82_n187), .A2(u5_mult_82_n70), 
        .ZN(u5_mult_82_FS_1_n200) );
  NAND4_X1 u5_mult_82_FS_1_U328 ( .A1(u5_mult_82_FS_1_n42), .A2(
        u5_mult_82_FS_1_n192), .A3(u5_mult_82_FS_1_n44), .A4(
        u5_mult_82_FS_1_n46), .ZN(u5_mult_82_FS_1_n188) );
  NOR2_X1 u5_mult_82_FS_1_U327 ( .A1(u5_mult_82_n186), .A2(u5_mult_82_n69), 
        .ZN(u5_mult_82_FS_1_n207) );
  NOR2_X1 u5_mult_82_FS_1_U326 ( .A1(u5_mult_82_n170), .A2(u5_mult_82_n68), 
        .ZN(u5_mult_82_FS_1_n214) );
  NAND2_X1 u5_mult_82_FS_1_U325 ( .A1(u5_mult_82_n169), .A2(u5_mult_82_n67), 
        .ZN(u5_mult_82_FS_1_n219) );
  NAND2_X1 u5_mult_82_FS_1_U324 ( .A1(u5_mult_82_n170), .A2(u5_mult_82_n68), 
        .ZN(u5_mult_82_FS_1_n216) );
  OAI21_X1 u5_mult_82_FS_1_U323 ( .B1(u5_mult_82_FS_1_n214), .B2(
        u5_mult_82_FS_1_n219), .A(u5_mult_82_FS_1_n216), .ZN(
        u5_mult_82_FS_1_n303) );
  NOR2_X1 u5_mult_82_FS_1_U322 ( .A1(u5_mult_82_n168), .A2(u5_mult_82_n66), 
        .ZN(u5_mult_82_FS_1_n209) );
  NAND2_X1 u5_mult_82_FS_1_U321 ( .A1(u5_mult_82_n168), .A2(u5_mult_82_n66), 
        .ZN(u5_mult_82_FS_1_n211) );
  AOI21_X1 u5_mult_82_FS_1_U320 ( .B1(u5_mult_82_FS_1_n303), .B2(
        u5_mult_82_FS_1_n51), .A(u5_mult_82_FS_1_n50), .ZN(
        u5_mult_82_FS_1_n302) );
  NAND2_X1 u5_mult_82_FS_1_U319 ( .A1(u5_mult_82_n186), .A2(u5_mult_82_n69), 
        .ZN(u5_mult_82_FS_1_n208) );
  OAI21_X1 u5_mult_82_FS_1_U318 ( .B1(u5_mult_82_FS_1_n207), .B2(
        u5_mult_82_FS_1_n302), .A(u5_mult_82_FS_1_n208), .ZN(
        u5_mult_82_FS_1_n203) );
  NOR2_X1 u5_mult_82_FS_1_U317 ( .A1(u5_mult_82_n162), .A2(u5_mult_82_n57), 
        .ZN(u5_mult_82_FS_1_n224) );
  NOR2_X1 u5_mult_82_FS_1_U316 ( .A1(u5_mult_82_n167), .A2(u5_mult_82_n65), 
        .ZN(u5_mult_82_FS_1_n228) );
  NOR2_X1 u5_mult_82_FS_1_U315 ( .A1(u5_mult_82_n161), .A2(u5_mult_82_n56), 
        .ZN(u5_mult_82_FS_1_n232) );
  NOR2_X1 u5_mult_82_FS_1_U314 ( .A1(u5_mult_82_n166), .A2(u5_mult_82_n64), 
        .ZN(u5_mult_82_FS_1_n236) );
  NOR2_X1 u5_mult_82_FS_1_U313 ( .A1(u5_mult_82_n165), .A2(u5_mult_82_n63), 
        .ZN(u5_mult_82_FS_1_n239) );
  OR2_X1 u5_mult_82_FS_1_U312 ( .A1(u5_mult_82_n160), .A2(u5_mult_82_n59), 
        .ZN(u5_mult_82_FS_1_n243) );
  NOR2_X1 u5_mult_82_FS_1_U311 ( .A1(u5_mult_82_n164), .A2(u5_mult_82_n62), 
        .ZN(u5_mult_82_FS_1_n247) );
  OR2_X1 u5_mult_82_FS_1_U310 ( .A1(u5_mult_82_n159), .A2(u5_mult_82_n58), 
        .ZN(u5_mult_82_FS_1_n251) );
  NOR2_X1 u5_mult_82_FS_1_U309 ( .A1(u5_mult_82_n163), .A2(u5_mult_82_n61), 
        .ZN(u5_mult_82_FS_1_n255) );
  NOR2_X1 u5_mult_82_FS_1_U308 ( .A1(u5_mult_82_n108), .A2(u5_mult_82_n7), 
        .ZN(u5_mult_82_FS_1_n260) );
  NOR2_X1 u5_mult_82_FS_1_U307 ( .A1(u5_mult_82_n106), .A2(u5_mult_82_n5), 
        .ZN(u5_mult_82_FS_1_n263) );
  NAND2_X1 u5_mult_82_FS_1_U306 ( .A1(u5_mult_82_n107), .A2(u5_mult_82_n6), 
        .ZN(u5_mult_82_FS_1_n264) );
  AND2_X1 u5_mult_82_FS_1_U305 ( .A1(u5_mult_82_n106), .A2(u5_mult_82_n5), 
        .ZN(u5_mult_82_FS_1_n262) );
  AOI21_X1 u5_mult_82_FS_1_U304 ( .B1(u5_mult_82_FS_1_n67), .B2(
        u5_mult_82_FS_1_n68), .A(u5_mult_82_FS_1_n262), .ZN(
        u5_mult_82_FS_1_n258) );
  NAND2_X1 u5_mult_82_FS_1_U303 ( .A1(u5_mult_82_n108), .A2(u5_mult_82_n7), 
        .ZN(u5_mult_82_FS_1_n259) );
  OAI21_X1 u5_mult_82_FS_1_U302 ( .B1(u5_mult_82_FS_1_n260), .B2(
        u5_mult_82_FS_1_n258), .A(u5_mult_82_FS_1_n259), .ZN(
        u5_mult_82_FS_1_n253) );
  NAND2_X1 u5_mult_82_FS_1_U301 ( .A1(u5_mult_82_n163), .A2(u5_mult_82_n61), 
        .ZN(u5_mult_82_FS_1_n256) );
  OAI21_X1 u5_mult_82_FS_1_U300 ( .B1(u5_mult_82_FS_1_n255), .B2(
        u5_mult_82_FS_1_n65), .A(u5_mult_82_FS_1_n256), .ZN(
        u5_mult_82_FS_1_n250) );
  NAND2_X1 u5_mult_82_FS_1_U299 ( .A1(u5_mult_82_n159), .A2(u5_mult_82_n58), 
        .ZN(u5_mult_82_FS_1_n252) );
  AOI21_X1 u5_mult_82_FS_1_U298 ( .B1(u5_mult_82_FS_1_n251), .B2(
        u5_mult_82_FS_1_n250), .A(u5_mult_82_FS_1_n63), .ZN(
        u5_mult_82_FS_1_n245) );
  NAND2_X1 u5_mult_82_FS_1_U297 ( .A1(u5_mult_82_n164), .A2(u5_mult_82_n62), 
        .ZN(u5_mult_82_FS_1_n248) );
  OAI21_X1 u5_mult_82_FS_1_U296 ( .B1(u5_mult_82_FS_1_n247), .B2(
        u5_mult_82_FS_1_n245), .A(u5_mult_82_FS_1_n248), .ZN(
        u5_mult_82_FS_1_n242) );
  NAND2_X1 u5_mult_82_FS_1_U295 ( .A1(u5_mult_82_n160), .A2(u5_mult_82_n59), 
        .ZN(u5_mult_82_FS_1_n244) );
  AOI21_X1 u5_mult_82_FS_1_U294 ( .B1(u5_mult_82_FS_1_n243), .B2(
        u5_mult_82_FS_1_n242), .A(u5_mult_82_FS_1_n61), .ZN(
        u5_mult_82_FS_1_n237) );
  NAND2_X1 u5_mult_82_FS_1_U293 ( .A1(u5_mult_82_n165), .A2(u5_mult_82_n63), 
        .ZN(u5_mult_82_FS_1_n240) );
  OAI21_X1 u5_mult_82_FS_1_U292 ( .B1(u5_mult_82_FS_1_n239), .B2(
        u5_mult_82_FS_1_n237), .A(u5_mult_82_FS_1_n240), .ZN(
        u5_mult_82_FS_1_n234) );
  NAND2_X1 u5_mult_82_FS_1_U291 ( .A1(u5_mult_82_n166), .A2(u5_mult_82_n64), 
        .ZN(u5_mult_82_FS_1_n235) );
  OAI21_X1 u5_mult_82_FS_1_U290 ( .B1(u5_mult_82_FS_1_n236), .B2(
        u5_mult_82_FS_1_n59), .A(u5_mult_82_FS_1_n235), .ZN(
        u5_mult_82_FS_1_n229) );
  AND2_X1 u5_mult_82_FS_1_U289 ( .A1(u5_mult_82_n161), .A2(u5_mult_82_n56), 
        .ZN(u5_mult_82_FS_1_n231) );
  AOI21_X1 u5_mult_82_FS_1_U288 ( .B1(u5_mult_82_FS_1_n57), .B2(
        u5_mult_82_FS_1_n229), .A(u5_mult_82_FS_1_n231), .ZN(
        u5_mult_82_FS_1_n226) );
  NAND2_X1 u5_mult_82_FS_1_U287 ( .A1(u5_mult_82_n167), .A2(u5_mult_82_n65), 
        .ZN(u5_mult_82_FS_1_n227) );
  OAI21_X1 u5_mult_82_FS_1_U286 ( .B1(u5_mult_82_FS_1_n228), .B2(
        u5_mult_82_FS_1_n226), .A(u5_mult_82_FS_1_n227), .ZN(
        u5_mult_82_FS_1_n221) );
  AND2_X1 u5_mult_82_FS_1_U285 ( .A1(u5_mult_82_n162), .A2(u5_mult_82_n57), 
        .ZN(u5_mult_82_FS_1_n223) );
  AOI21_X1 u5_mult_82_FS_1_U284 ( .B1(u5_mult_82_FS_1_n55), .B2(
        u5_mult_82_FS_1_n221), .A(u5_mult_82_FS_1_n223), .ZN(
        u5_mult_82_FS_1_n217) );
  NOR2_X1 u5_mult_82_FS_1_U283 ( .A1(u5_mult_82_n169), .A2(u5_mult_82_n67), 
        .ZN(u5_mult_82_FS_1_n218) );
  OR2_X1 u5_mult_82_FS_1_U282 ( .A1(u5_mult_82_FS_1_n217), .A2(
        u5_mult_82_FS_1_n218), .ZN(u5_mult_82_FS_1_n301) );
  NOR4_X1 u5_mult_82_FS_1_U281 ( .A1(u5_mult_82_FS_1_n207), .A2(
        u5_mult_82_FS_1_n209), .A3(u5_mult_82_FS_1_n301), .A4(
        u5_mult_82_FS_1_n214), .ZN(u5_mult_82_FS_1_n204) );
  NAND2_X1 u5_mult_82_FS_1_U280 ( .A1(u5_mult_82_n187), .A2(u5_mult_82_n70), 
        .ZN(u5_mult_82_FS_1_n201) );
  NAND2_X1 u5_mult_82_FS_1_U279 ( .A1(u5_mult_82_n188), .A2(u5_mult_82_n71), 
        .ZN(u5_mult_82_FS_1_n196) );
  OAI21_X1 u5_mult_82_FS_1_U278 ( .B1(u5_mult_82_FS_1_n195), .B2(
        u5_mult_82_FS_1_n201), .A(u5_mult_82_FS_1_n196), .ZN(
        u5_mult_82_FS_1_n300) );
  NAND2_X1 u5_mult_82_FS_1_U277 ( .A1(u5_mult_82_n172), .A2(u5_mult_82_n60), 
        .ZN(u5_mult_82_FS_1_n198) );
  AOI21_X1 u5_mult_82_FS_1_U276 ( .B1(u5_mult_82_FS_1_n300), .B2(
        u5_mult_82_FS_1_n192), .A(u5_mult_82_FS_1_n43), .ZN(
        u5_mult_82_FS_1_n299) );
  NAND2_X1 u5_mult_82_FS_1_U275 ( .A1(u5_mult_82_n189), .A2(u5_mult_82_n87), 
        .ZN(u5_mult_82_FS_1_n193) );
  OAI21_X1 u5_mult_82_FS_1_U274 ( .B1(u5_mult_82_FS_1_n298), .B2(
        u5_mult_82_FS_1_n299), .A(u5_mult_82_FS_1_n193), .ZN(
        u5_mult_82_FS_1_n297) );
  OAI221_X1 u5_mult_82_FS_1_U273 ( .B1(u5_mult_82_FS_1_n188), .B2(
        u5_mult_82_FS_1_n47), .C1(u5_mult_82_FS_1_n49), .C2(
        u5_mult_82_FS_1_n188), .A(u5_mult_82_FS_1_n41), .ZN(
        u5_mult_82_FS_1_n294) );
  NOR2_X1 u5_mult_82_FS_1_U272 ( .A1(u5_mult_82_n185), .A2(u5_mult_82_n86), 
        .ZN(u5_mult_82_FS_1_n177) );
  NOR2_X1 u5_mult_82_FS_1_U271 ( .A1(u5_mult_82_n174), .A2(u5_mult_82_n73), 
        .ZN(u5_mult_82_FS_1_n179) );
  NOR2_X1 u5_mult_82_FS_1_U270 ( .A1(u5_mult_82_n184), .A2(u5_mult_82_n85), 
        .ZN(u5_mult_82_FS_1_n180) );
  NOR2_X1 u5_mult_82_FS_1_U269 ( .A1(u5_mult_82_n183), .A2(u5_mult_82_n84), 
        .ZN(u5_mult_82_FS_1_n184) );
  NOR4_X1 u5_mult_82_FS_1_U268 ( .A1(u5_mult_82_FS_1_n177), .A2(
        u5_mult_82_FS_1_n179), .A3(u5_mult_82_FS_1_n180), .A4(
        u5_mult_82_FS_1_n184), .ZN(u5_mult_82_FS_1_n170) );
  NAND2_X1 u5_mult_82_FS_1_U267 ( .A1(u5_mult_82_n183), .A2(u5_mult_82_n84), 
        .ZN(u5_mult_82_FS_1_n186) );
  NAND2_X1 u5_mult_82_FS_1_U266 ( .A1(u5_mult_82_n184), .A2(u5_mult_82_n85), 
        .ZN(u5_mult_82_FS_1_n182) );
  OAI21_X1 u5_mult_82_FS_1_U265 ( .B1(u5_mult_82_FS_1_n180), .B2(
        u5_mult_82_FS_1_n186), .A(u5_mult_82_FS_1_n182), .ZN(
        u5_mult_82_FS_1_n296) );
  AND2_X1 u5_mult_82_FS_1_U264 ( .A1(u5_mult_82_n174), .A2(u5_mult_82_n73), 
        .ZN(u5_mult_82_FS_1_n175) );
  AOI21_X1 u5_mult_82_FS_1_U263 ( .B1(u5_mult_82_FS_1_n296), .B2(
        u5_mult_82_FS_1_n37), .A(u5_mult_82_FS_1_n175), .ZN(
        u5_mult_82_FS_1_n295) );
  NAND2_X1 u5_mult_82_FS_1_U262 ( .A1(u5_mult_82_n185), .A2(u5_mult_82_n86), 
        .ZN(u5_mult_82_FS_1_n176) );
  OAI21_X1 u5_mult_82_FS_1_U261 ( .B1(u5_mult_82_FS_1_n177), .B2(
        u5_mult_82_FS_1_n295), .A(u5_mult_82_FS_1_n176), .ZN(
        u5_mult_82_FS_1_n171) );
  AOI21_X1 u5_mult_82_FS_1_U260 ( .B1(u5_mult_82_FS_1_n294), .B2(
        u5_mult_82_FS_1_n170), .A(u5_mult_82_FS_1_n171), .ZN(
        u5_mult_82_FS_1_n293) );
  NOR2_X1 u5_mult_82_FS_1_U259 ( .A1(u5_mult_82_n182), .A2(u5_mult_82_n83), 
        .ZN(u5_mult_82_FS_1_n165) );
  NAND2_X1 u5_mult_82_FS_1_U258 ( .A1(u5_mult_82_n182), .A2(u5_mult_82_n83), 
        .ZN(u5_mult_82_FS_1_n167) );
  OAI21_X1 u5_mult_82_FS_1_U257 ( .B1(u5_mult_82_FS_1_n293), .B2(
        u5_mult_82_FS_1_n165), .A(u5_mult_82_FS_1_n167), .ZN(
        u5_mult_82_FS_1_n292) );
  AND2_X1 u5_mult_82_FS_1_U256 ( .A1(u5_mult_82_n175), .A2(u5_mult_82_n74), 
        .ZN(u5_mult_82_FS_1_n162) );
  AOI21_X1 u5_mult_82_FS_1_U255 ( .B1(u5_mult_82_FS_1_n34), .B2(
        u5_mult_82_FS_1_n292), .A(u5_mult_82_FS_1_n162), .ZN(
        u5_mult_82_FS_1_n291) );
  NOR2_X1 u5_mult_82_FS_1_U254 ( .A1(u5_mult_82_n181), .A2(u5_mult_82_n82), 
        .ZN(u5_mult_82_FS_1_n157) );
  NAND2_X1 u5_mult_82_FS_1_U253 ( .A1(u5_mult_82_n181), .A2(u5_mult_82_n82), 
        .ZN(u5_mult_82_FS_1_n159) );
  OAI21_X1 u5_mult_82_FS_1_U252 ( .B1(u5_mult_82_FS_1_n291), .B2(
        u5_mult_82_FS_1_n157), .A(u5_mult_82_FS_1_n159), .ZN(
        u5_mult_82_FS_1_n290) );
  AND2_X1 u5_mult_82_FS_1_U251 ( .A1(u5_mult_82_n176), .A2(u5_mult_82_n75), 
        .ZN(u5_mult_82_FS_1_n155) );
  AOI21_X1 u5_mult_82_FS_1_U250 ( .B1(u5_mult_82_FS_1_n32), .B2(
        u5_mult_82_FS_1_n290), .A(u5_mult_82_FS_1_n155), .ZN(
        u5_mult_82_FS_1_n149) );
  NAND2_X1 u5_mult_82_FS_1_U249 ( .A1(u5_mult_82_FS_1_n141), .A2(
        u5_mult_82_FS_1_n27), .ZN(u5_mult_82_FS_1_n288) );
  NOR4_X1 u5_mult_82_FS_1_U248 ( .A1(u5_mult_82_FS_1_n150), .A2(
        u5_mult_82_FS_1_n149), .A3(u5_mult_82_FS_1_n144), .A4(
        u5_mult_82_FS_1_n288), .ZN(u5_mult_82_FS_1_n137) );
  NAND2_X1 u5_mult_82_FS_1_U247 ( .A1(u5_mult_82_n193), .A2(u5_mult_82_n91), 
        .ZN(u5_mult_82_FS_1_n135) );
  NAND2_X1 u5_mult_82_FS_1_U246 ( .A1(u5_mult_82_n194), .A2(u5_mult_82_n92), 
        .ZN(u5_mult_82_FS_1_n131) );
  OAI21_X1 u5_mult_82_FS_1_U245 ( .B1(u5_mult_82_FS_1_n129), .B2(
        u5_mult_82_FS_1_n135), .A(u5_mult_82_FS_1_n131), .ZN(
        u5_mult_82_FS_1_n287) );
  AND2_X1 u5_mult_82_FS_1_U244 ( .A1(u5_mult_82_n177), .A2(u5_mult_82_n76), 
        .ZN(u5_mult_82_FS_1_n124) );
  AOI21_X1 u5_mult_82_FS_1_U243 ( .B1(u5_mult_82_FS_1_n287), .B2(
        u5_mult_82_FS_1_n23), .A(u5_mult_82_FS_1_n124), .ZN(
        u5_mult_82_FS_1_n286) );
  NAND2_X1 u5_mult_82_FS_1_U242 ( .A1(u5_mult_82_n195), .A2(u5_mult_82_n93), 
        .ZN(u5_mult_82_FS_1_n125) );
  OAI21_X1 u5_mult_82_FS_1_U241 ( .B1(u5_mult_82_FS_1_n126), .B2(
        u5_mult_82_FS_1_n286), .A(u5_mult_82_FS_1_n125), .ZN(
        u5_mult_82_FS_1_n120) );
  AOI221_X1 u5_mult_82_FS_1_U240 ( .B1(u5_mult_82_FS_1_n119), .B2(
        u5_mult_82_FS_1_n136), .C1(u5_mult_82_FS_1_n137), .C2(
        u5_mult_82_FS_1_n119), .A(u5_mult_82_FS_1_n120), .ZN(
        u5_mult_82_FS_1_n282) );
  NOR2_X1 u5_mult_82_FS_1_U239 ( .A1(u5_mult_82_n202), .A2(u5_mult_82_n81), 
        .ZN(u5_mult_82_FS_1_n105) );
  NOR2_X1 u5_mult_82_FS_1_U238 ( .A1(u5_mult_82_n180), .A2(u5_mult_82_n80), 
        .ZN(u5_mult_82_FS_1_n107) );
  NOR2_X1 u5_mult_82_FS_1_U237 ( .A1(u5_mult_82_n179), .A2(u5_mult_82_n79), 
        .ZN(u5_mult_82_FS_1_n112) );
  NOR2_X1 u5_mult_82_FS_1_U236 ( .A1(u5_mult_82_n178), .A2(u5_mult_82_n78), 
        .ZN(u5_mult_82_FS_1_n115) );
  OR4_X1 u5_mult_82_FS_1_U235 ( .A1(u5_mult_82_FS_1_n105), .A2(
        u5_mult_82_FS_1_n107), .A3(u5_mult_82_FS_1_n112), .A4(
        u5_mult_82_FS_1_n115), .ZN(u5_mult_82_FS_1_n102) );
  NAND2_X1 u5_mult_82_FS_1_U234 ( .A1(u5_mult_82_n178), .A2(u5_mult_82_n78), 
        .ZN(u5_mult_82_FS_1_n116) );
  NAND2_X1 u5_mult_82_FS_1_U233 ( .A1(u5_mult_82_n179), .A2(u5_mult_82_n79), 
        .ZN(u5_mult_82_FS_1_n114) );
  OAI21_X1 u5_mult_82_FS_1_U232 ( .B1(u5_mult_82_FS_1_n112), .B2(
        u5_mult_82_FS_1_n116), .A(u5_mult_82_FS_1_n114), .ZN(
        u5_mult_82_FS_1_n285) );
  NAND2_X1 u5_mult_82_FS_1_U231 ( .A1(u5_mult_82_n180), .A2(u5_mult_82_n80), 
        .ZN(u5_mult_82_FS_1_n109) );
  AOI21_X1 u5_mult_82_FS_1_U230 ( .B1(u5_mult_82_FS_1_n285), .B2(
        u5_mult_82_FS_1_n18), .A(u5_mult_82_FS_1_n17), .ZN(
        u5_mult_82_FS_1_n284) );
  NAND2_X1 u5_mult_82_FS_1_U229 ( .A1(u5_mult_82_n202), .A2(u5_mult_82_n81), 
        .ZN(u5_mult_82_FS_1_n106) );
  OAI21_X1 u5_mult_82_FS_1_U228 ( .B1(u5_mult_82_FS_1_n105), .B2(
        u5_mult_82_FS_1_n284), .A(u5_mult_82_FS_1_n106), .ZN(
        u5_mult_82_FS_1_n283) );
  OAI21_X1 u5_mult_82_FS_1_U227 ( .B1(u5_mult_82_FS_1_n282), .B2(
        u5_mult_82_FS_1_n102), .A(u5_mult_82_FS_1_n15), .ZN(
        u5_mult_82_FS_1_n281) );
  NOR2_X1 u5_mult_82_FS_1_U226 ( .A1(u5_mult_82_n199), .A2(u5_mult_82_n98), 
        .ZN(u5_mult_82_FS_1_n100) );
  AND2_X1 u5_mult_82_FS_1_U225 ( .A1(u5_mult_82_n199), .A2(u5_mult_82_n98), 
        .ZN(u5_mult_82_FS_1_n98) );
  AOI21_X1 u5_mult_82_FS_1_U224 ( .B1(u5_mult_82_FS_1_n281), .B2(
        u5_mult_82_FS_1_n14), .A(u5_mult_82_FS_1_n98), .ZN(
        u5_mult_82_FS_1_n280) );
  NAND2_X1 u5_mult_82_FS_1_U223 ( .A1(u5_mult_82_n203), .A2(u5_mult_82_n101), 
        .ZN(u5_mult_82_FS_1_n95) );
  OAI21_X1 u5_mult_82_FS_1_U222 ( .B1(u5_mult_82_FS_1_n93), .B2(
        u5_mult_82_FS_1_n280), .A(u5_mult_82_FS_1_n95), .ZN(
        u5_mult_82_FS_1_n279) );
  NOR2_X1 u5_mult_82_FS_1_U221 ( .A1(u5_mult_82_n198), .A2(u5_mult_82_n97), 
        .ZN(u5_mult_82_FS_1_n92) );
  AND2_X1 u5_mult_82_FS_1_U220 ( .A1(u5_mult_82_n198), .A2(u5_mult_82_n97), 
        .ZN(u5_mult_82_FS_1_n88) );
  AOI21_X1 u5_mult_82_FS_1_U219 ( .B1(u5_mult_82_FS_1_n279), .B2(
        u5_mult_82_FS_1_n12), .A(u5_mult_82_FS_1_n88), .ZN(
        u5_mult_82_FS_1_n278) );
  NAND2_X1 u5_mult_82_FS_1_U218 ( .A1(u5_mult_82_n204), .A2(u5_mult_82_n102), 
        .ZN(u5_mult_82_FS_1_n89) );
  OAI21_X1 u5_mult_82_FS_1_U217 ( .B1(u5_mult_82_FS_1_n90), .B2(
        u5_mult_82_FS_1_n278), .A(u5_mult_82_FS_1_n89), .ZN(
        u5_mult_82_FS_1_n82) );
  NOR2_X1 u5_mult_82_FS_1_U216 ( .A1(u5_mult_82_n201), .A2(u5_mult_82_n100), 
        .ZN(u5_mult_82_FS_1_n84) );
  NAND2_X1 u5_mult_82_FS_1_U215 ( .A1(u5_mult_82_n201), .A2(u5_mult_82_n100), 
        .ZN(u5_mult_82_FS_1_n83) );
  OAI21_X1 u5_mult_82_FS_1_U214 ( .B1(u5_mult_82_FS_1_n10), .B2(
        u5_mult_82_FS_1_n84), .A(u5_mult_82_FS_1_n83), .ZN(u5_mult_82_FS_1_n77) );
  AND2_X1 u5_mult_82_FS_1_U213 ( .A1(u5_mult_82_n200), .A2(u5_mult_82_n99), 
        .ZN(u5_mult_82_FS_1_n79) );
  AOI21_X1 u5_mult_82_FS_1_U212 ( .B1(u5_mult_82_FS_1_n8), .B2(
        u5_mult_82_FS_1_n77), .A(u5_mult_82_FS_1_n79), .ZN(u5_mult_82_FS_1_n74) );
  NAND2_X1 u5_mult_82_FS_1_U211 ( .A1(u5_mult_82_n205), .A2(u5_mult_82_n103), 
        .ZN(u5_mult_82_FS_1_n75) );
  OAI21_X1 u5_mult_82_FS_1_U210 ( .B1(u5_mult_82_FS_1_n76), .B2(
        u5_mult_82_FS_1_n74), .A(u5_mult_82_FS_1_n75), .ZN(u5_mult_82_FS_1_n69) );
  NOR2_X1 u5_mult_82_FS_1_U209 ( .A1(u5_mult_82_n197), .A2(u5_mult_82_n96), 
        .ZN(u5_mult_82_FS_1_n72) );
  AND2_X1 u5_mult_82_FS_1_U208 ( .A1(u5_mult_82_n197), .A2(u5_mult_82_n96), 
        .ZN(u5_mult_82_FS_1_n71) );
  AOI21_X1 u5_mult_82_FS_1_U207 ( .B1(u5_mult_82_FS_1_n69), .B2(
        u5_mult_82_FS_1_n6), .A(u5_mult_82_FS_1_n71), .ZN(u5_mult_82_FS_1_n275) );
  XOR2_X1 u5_mult_82_FS_1_U206 ( .A(u5_mult_82_FS_1_n277), .B(
        u5_mult_82_FS_1_n275), .Z(u5_N102) );
  OAI21_X1 u5_mult_82_FS_1_U205 ( .B1(u5_mult_82_FS_1_n274), .B2(
        u5_mult_82_FS_1_n275), .A(u5_mult_82_FS_1_n276), .ZN(
        u5_mult_82_FS_1_n270) );
  AND2_X1 u5_mult_82_FS_1_U204 ( .A1(u5_mult_82_n196), .A2(u5_mult_82_n95), 
        .ZN(u5_mult_82_FS_1_n271) );
  NOR2_X1 u5_mult_82_FS_1_U203 ( .A1(u5_mult_82_n196), .A2(u5_mult_82_n95), 
        .ZN(u5_mult_82_FS_1_n272) );
  NOR2_X1 u5_mult_82_FS_1_U202 ( .A1(u5_mult_82_FS_1_n271), .A2(
        u5_mult_82_FS_1_n272), .ZN(u5_mult_82_FS_1_n273) );
  XOR2_X1 u5_mult_82_FS_1_U201 ( .A(u5_mult_82_FS_1_n270), .B(
        u5_mult_82_FS_1_n273), .Z(u5_N103) );
  NOR2_X1 u5_mult_82_FS_1_U200 ( .A1(u5_mult_82_n209), .A2(u5_mult_82_n94), 
        .ZN(u5_mult_82_FS_1_n266) );
  NAND2_X1 u5_mult_82_FS_1_U199 ( .A1(u5_mult_82_n209), .A2(u5_mult_82_n94), 
        .ZN(u5_mult_82_FS_1_n268) );
  NAND2_X1 u5_mult_82_FS_1_U198 ( .A1(u5_mult_82_FS_1_n3), .A2(
        u5_mult_82_FS_1_n268), .ZN(u5_mult_82_FS_1_n269) );
  AOI21_X1 u5_mult_82_FS_1_U197 ( .B1(u5_mult_82_FS_1_n4), .B2(
        u5_mult_82_FS_1_n270), .A(u5_mult_82_FS_1_n271), .ZN(
        u5_mult_82_FS_1_n267) );
  XOR2_X1 u5_mult_82_FS_1_U196 ( .A(u5_mult_82_FS_1_n269), .B(
        u5_mult_82_FS_1_n267), .Z(u5_N104) );
  OAI21_X1 u5_mult_82_FS_1_U195 ( .B1(u5_mult_82_FS_1_n266), .B2(
        u5_mult_82_FS_1_n267), .A(u5_mult_82_FS_1_n268), .ZN(
        u5_mult_82_FS_1_n265) );
  XOR2_X1 u5_mult_82_FS_1_U194 ( .A(u5_mult_82_FS_1_n265), .B(u5_mult_82_n208), 
        .Z(u5_N105) );
  NOR2_X1 u5_mult_82_FS_1_U193 ( .A1(u5_mult_82_FS_1_n262), .A2(
        u5_mult_82_FS_1_n263), .ZN(u5_mult_82_FS_1_n261) );
  XOR2_X1 u5_mult_82_FS_1_U192 ( .A(u5_mult_82_FS_1_n68), .B(
        u5_mult_82_FS_1_n261), .Z(u5_N55) );
  NAND2_X1 u5_mult_82_FS_1_U191 ( .A1(u5_mult_82_FS_1_n66), .A2(
        u5_mult_82_FS_1_n259), .ZN(u5_mult_82_FS_1_n257) );
  XOR2_X1 u5_mult_82_FS_1_U190 ( .A(u5_mult_82_FS_1_n257), .B(
        u5_mult_82_FS_1_n258), .Z(u5_N56) );
  NOR2_X1 u5_mult_82_FS_1_U189 ( .A1(u5_mult_82_FS_1_n64), .A2(
        u5_mult_82_FS_1_n255), .ZN(u5_mult_82_FS_1_n254) );
  XOR2_X1 u5_mult_82_FS_1_U188 ( .A(u5_mult_82_FS_1_n253), .B(
        u5_mult_82_FS_1_n254), .Z(u5_N57) );
  NAND2_X1 u5_mult_82_FS_1_U187 ( .A1(u5_mult_82_FS_1_n251), .A2(
        u5_mult_82_FS_1_n252), .ZN(u5_mult_82_FS_1_n249) );
  XNOR2_X1 u5_mult_82_FS_1_U186 ( .A(u5_mult_82_FS_1_n249), .B(
        u5_mult_82_FS_1_n250), .ZN(u5_N58) );
  NOR2_X1 u5_mult_82_FS_1_U185 ( .A1(u5_mult_82_FS_1_n62), .A2(
        u5_mult_82_FS_1_n247), .ZN(u5_mult_82_FS_1_n246) );
  XNOR2_X1 u5_mult_82_FS_1_U184 ( .A(u5_mult_82_FS_1_n245), .B(
        u5_mult_82_FS_1_n246), .ZN(u5_N59) );
  NAND2_X1 u5_mult_82_FS_1_U183 ( .A1(u5_mult_82_FS_1_n243), .A2(
        u5_mult_82_FS_1_n244), .ZN(u5_mult_82_FS_1_n241) );
  XNOR2_X1 u5_mult_82_FS_1_U182 ( .A(u5_mult_82_FS_1_n241), .B(
        u5_mult_82_FS_1_n242), .ZN(u5_N60) );
  NOR2_X1 u5_mult_82_FS_1_U181 ( .A1(u5_mult_82_FS_1_n60), .A2(
        u5_mult_82_FS_1_n239), .ZN(u5_mult_82_FS_1_n238) );
  XNOR2_X1 u5_mult_82_FS_1_U180 ( .A(u5_mult_82_FS_1_n237), .B(
        u5_mult_82_FS_1_n238), .ZN(u5_N61) );
  NAND2_X1 u5_mult_82_FS_1_U179 ( .A1(u5_mult_82_FS_1_n58), .A2(
        u5_mult_82_FS_1_n235), .ZN(u5_mult_82_FS_1_n233) );
  XNOR2_X1 u5_mult_82_FS_1_U178 ( .A(u5_mult_82_FS_1_n233), .B(
        u5_mult_82_FS_1_n234), .ZN(u5_N62) );
  NOR2_X1 u5_mult_82_FS_1_U177 ( .A1(u5_mult_82_FS_1_n231), .A2(
        u5_mult_82_FS_1_n232), .ZN(u5_mult_82_FS_1_n230) );
  XOR2_X1 u5_mult_82_FS_1_U176 ( .A(u5_mult_82_FS_1_n229), .B(
        u5_mult_82_FS_1_n230), .Z(u5_N63) );
  NAND2_X1 u5_mult_82_FS_1_U175 ( .A1(u5_mult_82_FS_1_n56), .A2(
        u5_mult_82_FS_1_n227), .ZN(u5_mult_82_FS_1_n225) );
  XOR2_X1 u5_mult_82_FS_1_U174 ( .A(u5_mult_82_FS_1_n225), .B(
        u5_mult_82_FS_1_n226), .Z(u5_N64) );
  NOR2_X1 u5_mult_82_FS_1_U173 ( .A1(u5_mult_82_FS_1_n223), .A2(
        u5_mult_82_FS_1_n224), .ZN(u5_mult_82_FS_1_n222) );
  XOR2_X1 u5_mult_82_FS_1_U172 ( .A(u5_mult_82_FS_1_n221), .B(
        u5_mult_82_FS_1_n222), .Z(u5_N65) );
  NAND2_X1 u5_mult_82_FS_1_U171 ( .A1(u5_mult_82_FS_1_n54), .A2(
        u5_mult_82_FS_1_n219), .ZN(u5_mult_82_FS_1_n220) );
  XOR2_X1 u5_mult_82_FS_1_U170 ( .A(u5_mult_82_FS_1_n220), .B(
        u5_mult_82_FS_1_n217), .Z(u5_N66) );
  OAI21_X1 u5_mult_82_FS_1_U169 ( .B1(u5_mult_82_FS_1_n217), .B2(
        u5_mult_82_FS_1_n218), .A(u5_mult_82_FS_1_n219), .ZN(
        u5_mult_82_FS_1_n213) );
  NOR2_X1 u5_mult_82_FS_1_U168 ( .A1(u5_mult_82_FS_1_n52), .A2(
        u5_mult_82_FS_1_n214), .ZN(u5_mult_82_FS_1_n215) );
  XOR2_X1 u5_mult_82_FS_1_U167 ( .A(u5_mult_82_FS_1_n213), .B(
        u5_mult_82_FS_1_n215), .Z(u5_N67) );
  NAND2_X1 u5_mult_82_FS_1_U166 ( .A1(u5_mult_82_FS_1_n51), .A2(
        u5_mult_82_FS_1_n211), .ZN(u5_mult_82_FS_1_n212) );
  AOI21_X1 u5_mult_82_FS_1_U165 ( .B1(u5_mult_82_FS_1_n53), .B2(
        u5_mult_82_FS_1_n213), .A(u5_mult_82_FS_1_n52), .ZN(
        u5_mult_82_FS_1_n210) );
  XOR2_X1 u5_mult_82_FS_1_U164 ( .A(u5_mult_82_FS_1_n212), .B(
        u5_mult_82_FS_1_n210), .Z(u5_N68) );
  OAI21_X1 u5_mult_82_FS_1_U163 ( .B1(u5_mult_82_FS_1_n209), .B2(
        u5_mult_82_FS_1_n210), .A(u5_mult_82_FS_1_n211), .ZN(
        u5_mult_82_FS_1_n205) );
  NOR2_X1 u5_mult_82_FS_1_U162 ( .A1(u5_mult_82_FS_1_n48), .A2(
        u5_mult_82_FS_1_n207), .ZN(u5_mult_82_FS_1_n206) );
  XOR2_X1 u5_mult_82_FS_1_U161 ( .A(u5_mult_82_FS_1_n205), .B(
        u5_mult_82_FS_1_n206), .Z(u5_N69) );
  NAND2_X1 u5_mult_82_FS_1_U160 ( .A1(u5_mult_82_FS_1_n46), .A2(
        u5_mult_82_FS_1_n201), .ZN(u5_mult_82_FS_1_n202) );
  NOR2_X1 u5_mult_82_FS_1_U159 ( .A1(u5_mult_82_FS_1_n203), .A2(
        u5_mult_82_FS_1_n204), .ZN(u5_mult_82_FS_1_n187) );
  XOR2_X1 u5_mult_82_FS_1_U158 ( .A(u5_mult_82_FS_1_n202), .B(
        u5_mult_82_FS_1_n187), .Z(u5_N70) );
  NAND2_X1 u5_mult_82_FS_1_U157 ( .A1(u5_mult_82_FS_1_n44), .A2(
        u5_mult_82_FS_1_n196), .ZN(u5_mult_82_FS_1_n199) );
  OAI21_X1 u5_mult_82_FS_1_U156 ( .B1(u5_mult_82_FS_1_n200), .B2(
        u5_mult_82_FS_1_n187), .A(u5_mult_82_FS_1_n201), .ZN(
        u5_mult_82_FS_1_n197) );
  XNOR2_X1 u5_mult_82_FS_1_U155 ( .A(u5_mult_82_FS_1_n199), .B(
        u5_mult_82_FS_1_n197), .ZN(u5_N71) );
  NAND2_X1 u5_mult_82_FS_1_U154 ( .A1(u5_mult_82_FS_1_n192), .A2(
        u5_mult_82_FS_1_n198), .ZN(u5_mult_82_FS_1_n194) );
  OAI21_X1 u5_mult_82_FS_1_U153 ( .B1(u5_mult_82_FS_1_n195), .B2(
        u5_mult_82_FS_1_n45), .A(u5_mult_82_FS_1_n196), .ZN(
        u5_mult_82_FS_1_n191) );
  XNOR2_X1 u5_mult_82_FS_1_U152 ( .A(u5_mult_82_FS_1_n194), .B(
        u5_mult_82_FS_1_n191), .ZN(u5_N72) );
  NAND2_X1 u5_mult_82_FS_1_U151 ( .A1(u5_mult_82_FS_1_n42), .A2(
        u5_mult_82_FS_1_n193), .ZN(u5_mult_82_FS_1_n189) );
  AOI21_X1 u5_mult_82_FS_1_U150 ( .B1(u5_mult_82_FS_1_n191), .B2(
        u5_mult_82_FS_1_n192), .A(u5_mult_82_FS_1_n43), .ZN(
        u5_mult_82_FS_1_n190) );
  XOR2_X1 u5_mult_82_FS_1_U149 ( .A(u5_mult_82_FS_1_n189), .B(
        u5_mult_82_FS_1_n190), .Z(u5_N73) );
  OAI21_X1 u5_mult_82_FS_1_U148 ( .B1(u5_mult_82_FS_1_n187), .B2(
        u5_mult_82_FS_1_n188), .A(u5_mult_82_FS_1_n41), .ZN(
        u5_mult_82_FS_1_n169) );
  NOR2_X1 u5_mult_82_FS_1_U147 ( .A1(u5_mult_82_FS_1_n39), .A2(
        u5_mult_82_FS_1_n184), .ZN(u5_mult_82_FS_1_n185) );
  XOR2_X1 u5_mult_82_FS_1_U146 ( .A(u5_mult_82_FS_1_n169), .B(
        u5_mult_82_FS_1_n185), .Z(u5_N74) );
  NAND2_X1 u5_mult_82_FS_1_U145 ( .A1(u5_mult_82_FS_1_n38), .A2(
        u5_mult_82_FS_1_n182), .ZN(u5_mult_82_FS_1_n183) );
  AOI21_X1 u5_mult_82_FS_1_U144 ( .B1(u5_mult_82_FS_1_n40), .B2(
        u5_mult_82_FS_1_n169), .A(u5_mult_82_FS_1_n39), .ZN(
        u5_mult_82_FS_1_n181) );
  XOR2_X1 u5_mult_82_FS_1_U143 ( .A(u5_mult_82_FS_1_n183), .B(
        u5_mult_82_FS_1_n181), .Z(u5_N75) );
  OAI21_X1 u5_mult_82_FS_1_U142 ( .B1(u5_mult_82_FS_1_n180), .B2(
        u5_mult_82_FS_1_n181), .A(u5_mult_82_FS_1_n182), .ZN(
        u5_mult_82_FS_1_n174) );
  NOR2_X1 u5_mult_82_FS_1_U141 ( .A1(u5_mult_82_FS_1_n175), .A2(
        u5_mult_82_FS_1_n179), .ZN(u5_mult_82_FS_1_n178) );
  XOR2_X1 u5_mult_82_FS_1_U140 ( .A(u5_mult_82_FS_1_n174), .B(
        u5_mult_82_FS_1_n178), .Z(u5_N76) );
  NAND2_X1 u5_mult_82_FS_1_U139 ( .A1(u5_mult_82_FS_1_n36), .A2(
        u5_mult_82_FS_1_n176), .ZN(u5_mult_82_FS_1_n172) );
  AOI21_X1 u5_mult_82_FS_1_U138 ( .B1(u5_mult_82_FS_1_n174), .B2(
        u5_mult_82_FS_1_n37), .A(u5_mult_82_FS_1_n175), .ZN(
        u5_mult_82_FS_1_n173) );
  XOR2_X1 u5_mult_82_FS_1_U137 ( .A(u5_mult_82_FS_1_n172), .B(
        u5_mult_82_FS_1_n173), .Z(u5_N77) );
  NAND2_X1 u5_mult_82_FS_1_U136 ( .A1(u5_mult_82_FS_1_n35), .A2(
        u5_mult_82_FS_1_n167), .ZN(u5_mult_82_FS_1_n168) );
  AOI21_X1 u5_mult_82_FS_1_U135 ( .B1(u5_mult_82_FS_1_n169), .B2(
        u5_mult_82_FS_1_n170), .A(u5_mult_82_FS_1_n171), .ZN(
        u5_mult_82_FS_1_n166) );
  XOR2_X1 u5_mult_82_FS_1_U134 ( .A(u5_mult_82_FS_1_n168), .B(
        u5_mult_82_FS_1_n166), .Z(u5_N78) );
  OAI21_X1 u5_mult_82_FS_1_U133 ( .B1(u5_mult_82_FS_1_n165), .B2(
        u5_mult_82_FS_1_n166), .A(u5_mult_82_FS_1_n167), .ZN(
        u5_mult_82_FS_1_n161) );
  NOR2_X1 u5_mult_82_FS_1_U132 ( .A1(u5_mult_82_FS_1_n162), .A2(
        u5_mult_82_FS_1_n164), .ZN(u5_mult_82_FS_1_n163) );
  XOR2_X1 u5_mult_82_FS_1_U131 ( .A(u5_mult_82_FS_1_n161), .B(
        u5_mult_82_FS_1_n163), .Z(u5_N79) );
  NAND2_X1 u5_mult_82_FS_1_U130 ( .A1(u5_mult_82_FS_1_n33), .A2(
        u5_mult_82_FS_1_n159), .ZN(u5_mult_82_FS_1_n160) );
  AOI21_X1 u5_mult_82_FS_1_U129 ( .B1(u5_mult_82_FS_1_n34), .B2(
        u5_mult_82_FS_1_n161), .A(u5_mult_82_FS_1_n162), .ZN(
        u5_mult_82_FS_1_n158) );
  XOR2_X1 u5_mult_82_FS_1_U128 ( .A(u5_mult_82_FS_1_n160), .B(
        u5_mult_82_FS_1_n158), .Z(u5_N80) );
  OAI21_X1 u5_mult_82_FS_1_U127 ( .B1(u5_mult_82_FS_1_n157), .B2(
        u5_mult_82_FS_1_n158), .A(u5_mult_82_FS_1_n159), .ZN(
        u5_mult_82_FS_1_n153) );
  NOR2_X1 u5_mult_82_FS_1_U126 ( .A1(u5_mult_82_FS_1_n155), .A2(
        u5_mult_82_FS_1_n156), .ZN(u5_mult_82_FS_1_n154) );
  XOR2_X1 u5_mult_82_FS_1_U125 ( .A(u5_mult_82_FS_1_n153), .B(
        u5_mult_82_FS_1_n154), .Z(u5_N81) );
  NOR2_X1 u5_mult_82_FS_1_U124 ( .A1(u5_mult_82_FS_1_n31), .A2(
        u5_mult_82_FS_1_n150), .ZN(u5_mult_82_FS_1_n152) );
  XNOR2_X1 u5_mult_82_FS_1_U123 ( .A(u5_mult_82_FS_1_n149), .B(
        u5_mult_82_FS_1_n152), .ZN(u5_N82) );
  NAND2_X1 u5_mult_82_FS_1_U122 ( .A1(u5_mult_82_FS_1_n29), .A2(
        u5_mult_82_FS_1_n145), .ZN(u5_mult_82_FS_1_n147) );
  OAI21_X1 u5_mult_82_FS_1_U121 ( .B1(u5_mult_82_FS_1_n149), .B2(
        u5_mult_82_FS_1_n150), .A(u5_mult_82_FS_1_n151), .ZN(
        u5_mult_82_FS_1_n148) );
  XOR2_X1 u5_mult_82_FS_1_U120 ( .A(u5_mult_82_FS_1_n147), .B(
        u5_mult_82_FS_1_n30), .Z(u5_N83) );
  NAND2_X1 u5_mult_82_FS_1_U119 ( .A1(u5_mult_82_FS_1_n141), .A2(
        u5_mult_82_FS_1_n146), .ZN(u5_mult_82_FS_1_n143) );
  OAI21_X1 u5_mult_82_FS_1_U118 ( .B1(u5_mult_82_FS_1_n144), .B2(
        u5_mult_82_FS_1_n30), .A(u5_mult_82_FS_1_n145), .ZN(
        u5_mult_82_FS_1_n140) );
  XNOR2_X1 u5_mult_82_FS_1_U117 ( .A(u5_mult_82_FS_1_n143), .B(
        u5_mult_82_FS_1_n140), .ZN(u5_N84) );
  NAND2_X1 u5_mult_82_FS_1_U116 ( .A1(u5_mult_82_FS_1_n27), .A2(
        u5_mult_82_FS_1_n142), .ZN(u5_mult_82_FS_1_n138) );
  AOI21_X1 u5_mult_82_FS_1_U115 ( .B1(u5_mult_82_FS_1_n140), .B2(
        u5_mult_82_FS_1_n141), .A(u5_mult_82_FS_1_n28), .ZN(
        u5_mult_82_FS_1_n139) );
  XOR2_X1 u5_mult_82_FS_1_U114 ( .A(u5_mult_82_FS_1_n138), .B(
        u5_mult_82_FS_1_n139), .Z(u5_N85) );
  OR2_X1 u5_mult_82_FS_1_U113 ( .A1(u5_mult_82_FS_1_n136), .A2(
        u5_mult_82_FS_1_n137), .ZN(u5_mult_82_FS_1_n118) );
  NOR2_X1 u5_mult_82_FS_1_U112 ( .A1(u5_mult_82_FS_1_n25), .A2(
        u5_mult_82_FS_1_n133), .ZN(u5_mult_82_FS_1_n134) );
  XOR2_X1 u5_mult_82_FS_1_U111 ( .A(u5_mult_82_FS_1_n118), .B(
        u5_mult_82_FS_1_n134), .Z(u5_N86) );
  NAND2_X1 u5_mult_82_FS_1_U110 ( .A1(u5_mult_82_FS_1_n24), .A2(
        u5_mult_82_FS_1_n131), .ZN(u5_mult_82_FS_1_n132) );
  AOI21_X1 u5_mult_82_FS_1_U109 ( .B1(u5_mult_82_FS_1_n26), .B2(
        u5_mult_82_FS_1_n118), .A(u5_mult_82_FS_1_n25), .ZN(
        u5_mult_82_FS_1_n130) );
  XOR2_X1 u5_mult_82_FS_1_U108 ( .A(u5_mult_82_FS_1_n132), .B(
        u5_mult_82_FS_1_n130), .Z(u5_N87) );
  OAI21_X1 u5_mult_82_FS_1_U107 ( .B1(u5_mult_82_FS_1_n129), .B2(
        u5_mult_82_FS_1_n130), .A(u5_mult_82_FS_1_n131), .ZN(
        u5_mult_82_FS_1_n123) );
  NOR2_X1 u5_mult_82_FS_1_U106 ( .A1(u5_mult_82_FS_1_n124), .A2(
        u5_mult_82_FS_1_n128), .ZN(u5_mult_82_FS_1_n127) );
  XOR2_X1 u5_mult_82_FS_1_U105 ( .A(u5_mult_82_FS_1_n123), .B(
        u5_mult_82_FS_1_n127), .Z(u5_N88) );
  NAND2_X1 u5_mult_82_FS_1_U104 ( .A1(u5_mult_82_FS_1_n22), .A2(
        u5_mult_82_FS_1_n125), .ZN(u5_mult_82_FS_1_n121) );
  AOI21_X1 u5_mult_82_FS_1_U103 ( .B1(u5_mult_82_FS_1_n123), .B2(
        u5_mult_82_FS_1_n23), .A(u5_mult_82_FS_1_n124), .ZN(
        u5_mult_82_FS_1_n122) );
  XOR2_X1 u5_mult_82_FS_1_U102 ( .A(u5_mult_82_FS_1_n121), .B(
        u5_mult_82_FS_1_n122), .Z(u5_N89) );
  NAND2_X1 u5_mult_82_FS_1_U101 ( .A1(u5_mult_82_FS_1_n21), .A2(
        u5_mult_82_FS_1_n116), .ZN(u5_mult_82_FS_1_n117) );
  AOI21_X1 u5_mult_82_FS_1_U100 ( .B1(u5_mult_82_FS_1_n118), .B2(
        u5_mult_82_FS_1_n119), .A(u5_mult_82_FS_1_n120), .ZN(
        u5_mult_82_FS_1_n101) );
  XOR2_X1 u5_mult_82_FS_1_U99 ( .A(u5_mult_82_FS_1_n117), .B(
        u5_mult_82_FS_1_n101), .Z(u5_N90) );
  OAI21_X1 u5_mult_82_FS_1_U98 ( .B1(u5_mult_82_FS_1_n115), .B2(
        u5_mult_82_FS_1_n101), .A(u5_mult_82_FS_1_n116), .ZN(
        u5_mult_82_FS_1_n111) );
  NOR2_X1 u5_mult_82_FS_1_U97 ( .A1(u5_mult_82_FS_1_n19), .A2(
        u5_mult_82_FS_1_n112), .ZN(u5_mult_82_FS_1_n113) );
  XOR2_X1 u5_mult_82_FS_1_U96 ( .A(u5_mult_82_FS_1_n111), .B(
        u5_mult_82_FS_1_n113), .Z(u5_N91) );
  NAND2_X1 u5_mult_82_FS_1_U95 ( .A1(u5_mult_82_FS_1_n18), .A2(
        u5_mult_82_FS_1_n109), .ZN(u5_mult_82_FS_1_n110) );
  AOI21_X1 u5_mult_82_FS_1_U94 ( .B1(u5_mult_82_FS_1_n20), .B2(
        u5_mult_82_FS_1_n111), .A(u5_mult_82_FS_1_n19), .ZN(
        u5_mult_82_FS_1_n108) );
  XOR2_X1 u5_mult_82_FS_1_U93 ( .A(u5_mult_82_FS_1_n110), .B(
        u5_mult_82_FS_1_n108), .Z(u5_N92) );
  OAI21_X1 u5_mult_82_FS_1_U92 ( .B1(u5_mult_82_FS_1_n107), .B2(
        u5_mult_82_FS_1_n108), .A(u5_mult_82_FS_1_n109), .ZN(
        u5_mult_82_FS_1_n103) );
  NOR2_X1 u5_mult_82_FS_1_U91 ( .A1(u5_mult_82_FS_1_n16), .A2(
        u5_mult_82_FS_1_n105), .ZN(u5_mult_82_FS_1_n104) );
  XOR2_X1 u5_mult_82_FS_1_U90 ( .A(u5_mult_82_FS_1_n103), .B(
        u5_mult_82_FS_1_n104), .Z(u5_N93) );
  OAI21_X1 u5_mult_82_FS_1_U89 ( .B1(u5_mult_82_FS_1_n101), .B2(
        u5_mult_82_FS_1_n102), .A(u5_mult_82_FS_1_n15), .ZN(
        u5_mult_82_FS_1_n97) );
  NOR2_X1 u5_mult_82_FS_1_U88 ( .A1(u5_mult_82_FS_1_n98), .A2(
        u5_mult_82_FS_1_n100), .ZN(u5_mult_82_FS_1_n99) );
  XOR2_X1 u5_mult_82_FS_1_U87 ( .A(u5_mult_82_FS_1_n97), .B(
        u5_mult_82_FS_1_n99), .Z(u5_N94) );
  NAND2_X1 u5_mult_82_FS_1_U86 ( .A1(u5_mult_82_FS_1_n13), .A2(
        u5_mult_82_FS_1_n95), .ZN(u5_mult_82_FS_1_n96) );
  AOI21_X1 u5_mult_82_FS_1_U85 ( .B1(u5_mult_82_FS_1_n14), .B2(
        u5_mult_82_FS_1_n97), .A(u5_mult_82_FS_1_n98), .ZN(u5_mult_82_FS_1_n94) );
  XOR2_X1 u5_mult_82_FS_1_U84 ( .A(u5_mult_82_FS_1_n96), .B(
        u5_mult_82_FS_1_n94), .Z(u5_N95) );
  OAI21_X1 u5_mult_82_FS_1_U83 ( .B1(u5_mult_82_FS_1_n93), .B2(
        u5_mult_82_FS_1_n94), .A(u5_mult_82_FS_1_n95), .ZN(u5_mult_82_FS_1_n87) );
  NOR2_X1 u5_mult_82_FS_1_U82 ( .A1(u5_mult_82_FS_1_n88), .A2(
        u5_mult_82_FS_1_n92), .ZN(u5_mult_82_FS_1_n91) );
  XOR2_X1 u5_mult_82_FS_1_U81 ( .A(u5_mult_82_FS_1_n87), .B(
        u5_mult_82_FS_1_n91), .Z(u5_N96) );
  NAND2_X1 u5_mult_82_FS_1_U80 ( .A1(u5_mult_82_FS_1_n11), .A2(
        u5_mult_82_FS_1_n89), .ZN(u5_mult_82_FS_1_n85) );
  AOI21_X1 u5_mult_82_FS_1_U79 ( .B1(u5_mult_82_FS_1_n87), .B2(
        u5_mult_82_FS_1_n12), .A(u5_mult_82_FS_1_n88), .ZN(u5_mult_82_FS_1_n86) );
  XOR2_X1 u5_mult_82_FS_1_U78 ( .A(u5_mult_82_FS_1_n85), .B(
        u5_mult_82_FS_1_n86), .Z(u5_N97) );
  NAND2_X1 u5_mult_82_FS_1_U77 ( .A1(u5_mult_82_FS_1_n9), .A2(
        u5_mult_82_FS_1_n83), .ZN(u5_mult_82_FS_1_n81) );
  XNOR2_X1 u5_mult_82_FS_1_U76 ( .A(u5_mult_82_FS_1_n81), .B(
        u5_mult_82_FS_1_n82), .ZN(u5_N98) );
  NOR2_X1 u5_mult_82_FS_1_U75 ( .A1(u5_mult_82_FS_1_n79), .A2(
        u5_mult_82_FS_1_n80), .ZN(u5_mult_82_FS_1_n78) );
  XOR2_X1 u5_mult_82_FS_1_U74 ( .A(u5_mult_82_FS_1_n77), .B(
        u5_mult_82_FS_1_n78), .Z(u5_N99) );
  NAND2_X1 u5_mult_82_FS_1_U73 ( .A1(u5_mult_82_FS_1_n7), .A2(
        u5_mult_82_FS_1_n75), .ZN(u5_mult_82_FS_1_n73) );
  XOR2_X1 u5_mult_82_FS_1_U72 ( .A(u5_mult_82_FS_1_n73), .B(
        u5_mult_82_FS_1_n74), .Z(u5_N100) );
  NOR2_X1 u5_mult_82_FS_1_U71 ( .A1(u5_mult_82_FS_1_n71), .A2(
        u5_mult_82_FS_1_n72), .ZN(u5_mult_82_FS_1_n70) );
  XOR2_X1 u5_mult_82_FS_1_U70 ( .A(u5_mult_82_FS_1_n69), .B(
        u5_mult_82_FS_1_n70), .Z(u5_N101) );
  INV_X4 u5_mult_82_FS_1_U69 ( .A(u5_mult_82_FS_1_n264), .ZN(
        u5_mult_82_FS_1_n68) );
  INV_X4 u5_mult_82_FS_1_U68 ( .A(u5_mult_82_FS_1_n263), .ZN(
        u5_mult_82_FS_1_n67) );
  INV_X4 u5_mult_82_FS_1_U67 ( .A(u5_mult_82_FS_1_n260), .ZN(
        u5_mult_82_FS_1_n66) );
  INV_X4 u5_mult_82_FS_1_U66 ( .A(u5_mult_82_FS_1_n253), .ZN(
        u5_mult_82_FS_1_n65) );
  INV_X4 u5_mult_82_FS_1_U65 ( .A(u5_mult_82_FS_1_n256), .ZN(
        u5_mult_82_FS_1_n64) );
  INV_X4 u5_mult_82_FS_1_U64 ( .A(u5_mult_82_FS_1_n252), .ZN(
        u5_mult_82_FS_1_n63) );
  INV_X4 u5_mult_82_FS_1_U63 ( .A(u5_mult_82_FS_1_n248), .ZN(
        u5_mult_82_FS_1_n62) );
  INV_X4 u5_mult_82_FS_1_U62 ( .A(u5_mult_82_FS_1_n244), .ZN(
        u5_mult_82_FS_1_n61) );
  INV_X4 u5_mult_82_FS_1_U61 ( .A(u5_mult_82_FS_1_n240), .ZN(
        u5_mult_82_FS_1_n60) );
  INV_X4 u5_mult_82_FS_1_U60 ( .A(u5_mult_82_FS_1_n234), .ZN(
        u5_mult_82_FS_1_n59) );
  INV_X4 u5_mult_82_FS_1_U59 ( .A(u5_mult_82_FS_1_n236), .ZN(
        u5_mult_82_FS_1_n58) );
  INV_X4 u5_mult_82_FS_1_U58 ( .A(u5_mult_82_FS_1_n232), .ZN(
        u5_mult_82_FS_1_n57) );
  INV_X4 u5_mult_82_FS_1_U57 ( .A(u5_mult_82_FS_1_n228), .ZN(
        u5_mult_82_FS_1_n56) );
  INV_X4 u5_mult_82_FS_1_U56 ( .A(u5_mult_82_FS_1_n224), .ZN(
        u5_mult_82_FS_1_n55) );
  INV_X4 u5_mult_82_FS_1_U55 ( .A(u5_mult_82_FS_1_n218), .ZN(
        u5_mult_82_FS_1_n54) );
  INV_X4 u5_mult_82_FS_1_U54 ( .A(u5_mult_82_FS_1_n214), .ZN(
        u5_mult_82_FS_1_n53) );
  INV_X4 u5_mult_82_FS_1_U53 ( .A(u5_mult_82_FS_1_n216), .ZN(
        u5_mult_82_FS_1_n52) );
  INV_X4 u5_mult_82_FS_1_U52 ( .A(u5_mult_82_FS_1_n209), .ZN(
        u5_mult_82_FS_1_n51) );
  INV_X4 u5_mult_82_FS_1_U51 ( .A(u5_mult_82_FS_1_n211), .ZN(
        u5_mult_82_FS_1_n50) );
  INV_X4 u5_mult_82_FS_1_U50 ( .A(u5_mult_82_FS_1_n204), .ZN(
        u5_mult_82_FS_1_n49) );
  INV_X4 u5_mult_82_FS_1_U49 ( .A(u5_mult_82_FS_1_n208), .ZN(
        u5_mult_82_FS_1_n48) );
  INV_X4 u5_mult_82_FS_1_U48 ( .A(u5_mult_82_FS_1_n203), .ZN(
        u5_mult_82_FS_1_n47) );
  INV_X4 u5_mult_82_FS_1_U47 ( .A(u5_mult_82_FS_1_n200), .ZN(
        u5_mult_82_FS_1_n46) );
  INV_X4 u5_mult_82_FS_1_U46 ( .A(u5_mult_82_FS_1_n197), .ZN(
        u5_mult_82_FS_1_n45) );
  INV_X4 u5_mult_82_FS_1_U45 ( .A(u5_mult_82_FS_1_n195), .ZN(
        u5_mult_82_FS_1_n44) );
  INV_X4 u5_mult_82_FS_1_U44 ( .A(u5_mult_82_FS_1_n198), .ZN(
        u5_mult_82_FS_1_n43) );
  INV_X4 u5_mult_82_FS_1_U43 ( .A(u5_mult_82_FS_1_n298), .ZN(
        u5_mult_82_FS_1_n42) );
  INV_X4 u5_mult_82_FS_1_U42 ( .A(u5_mult_82_FS_1_n297), .ZN(
        u5_mult_82_FS_1_n41) );
  INV_X4 u5_mult_82_FS_1_U41 ( .A(u5_mult_82_FS_1_n184), .ZN(
        u5_mult_82_FS_1_n40) );
  INV_X4 u5_mult_82_FS_1_U40 ( .A(u5_mult_82_FS_1_n186), .ZN(
        u5_mult_82_FS_1_n39) );
  INV_X4 u5_mult_82_FS_1_U39 ( .A(u5_mult_82_FS_1_n180), .ZN(
        u5_mult_82_FS_1_n38) );
  INV_X4 u5_mult_82_FS_1_U38 ( .A(u5_mult_82_FS_1_n179), .ZN(
        u5_mult_82_FS_1_n37) );
  INV_X4 u5_mult_82_FS_1_U37 ( .A(u5_mult_82_FS_1_n177), .ZN(
        u5_mult_82_FS_1_n36) );
  INV_X4 u5_mult_82_FS_1_U36 ( .A(u5_mult_82_FS_1_n165), .ZN(
        u5_mult_82_FS_1_n35) );
  INV_X4 u5_mult_82_FS_1_U35 ( .A(u5_mult_82_FS_1_n164), .ZN(
        u5_mult_82_FS_1_n34) );
  INV_X4 u5_mult_82_FS_1_U34 ( .A(u5_mult_82_FS_1_n157), .ZN(
        u5_mult_82_FS_1_n33) );
  INV_X4 u5_mult_82_FS_1_U33 ( .A(u5_mult_82_FS_1_n156), .ZN(
        u5_mult_82_FS_1_n32) );
  INV_X4 u5_mult_82_FS_1_U32 ( .A(u5_mult_82_FS_1_n151), .ZN(
        u5_mult_82_FS_1_n31) );
  INV_X4 u5_mult_82_FS_1_U31 ( .A(u5_mult_82_FS_1_n148), .ZN(
        u5_mult_82_FS_1_n30) );
  INV_X4 u5_mult_82_FS_1_U30 ( .A(u5_mult_82_FS_1_n144), .ZN(
        u5_mult_82_FS_1_n29) );
  INV_X4 u5_mult_82_FS_1_U29 ( .A(u5_mult_82_FS_1_n146), .ZN(
        u5_mult_82_FS_1_n28) );
  INV_X4 u5_mult_82_FS_1_U28 ( .A(u5_mult_82_FS_1_n289), .ZN(
        u5_mult_82_FS_1_n27) );
  INV_X4 u5_mult_82_FS_1_U27 ( .A(u5_mult_82_FS_1_n133), .ZN(
        u5_mult_82_FS_1_n26) );
  INV_X4 u5_mult_82_FS_1_U26 ( .A(u5_mult_82_FS_1_n135), .ZN(
        u5_mult_82_FS_1_n25) );
  INV_X4 u5_mult_82_FS_1_U25 ( .A(u5_mult_82_FS_1_n129), .ZN(
        u5_mult_82_FS_1_n24) );
  INV_X4 u5_mult_82_FS_1_U24 ( .A(u5_mult_82_FS_1_n128), .ZN(
        u5_mult_82_FS_1_n23) );
  INV_X4 u5_mult_82_FS_1_U23 ( .A(u5_mult_82_FS_1_n126), .ZN(
        u5_mult_82_FS_1_n22) );
  INV_X4 u5_mult_82_FS_1_U22 ( .A(u5_mult_82_FS_1_n115), .ZN(
        u5_mult_82_FS_1_n21) );
  INV_X4 u5_mult_82_FS_1_U21 ( .A(u5_mult_82_FS_1_n112), .ZN(
        u5_mult_82_FS_1_n20) );
  INV_X4 u5_mult_82_FS_1_U20 ( .A(u5_mult_82_FS_1_n114), .ZN(
        u5_mult_82_FS_1_n19) );
  INV_X4 u5_mult_82_FS_1_U19 ( .A(u5_mult_82_FS_1_n107), .ZN(
        u5_mult_82_FS_1_n18) );
  INV_X4 u5_mult_82_FS_1_U18 ( .A(u5_mult_82_FS_1_n109), .ZN(
        u5_mult_82_FS_1_n17) );
  INV_X4 u5_mult_82_FS_1_U17 ( .A(u5_mult_82_FS_1_n106), .ZN(
        u5_mult_82_FS_1_n16) );
  INV_X4 u5_mult_82_FS_1_U16 ( .A(u5_mult_82_FS_1_n283), .ZN(
        u5_mult_82_FS_1_n15) );
  INV_X4 u5_mult_82_FS_1_U15 ( .A(u5_mult_82_FS_1_n100), .ZN(
        u5_mult_82_FS_1_n14) );
  INV_X4 u5_mult_82_FS_1_U14 ( .A(u5_mult_82_FS_1_n93), .ZN(
        u5_mult_82_FS_1_n13) );
  INV_X4 u5_mult_82_FS_1_U13 ( .A(u5_mult_82_FS_1_n92), .ZN(
        u5_mult_82_FS_1_n12) );
  INV_X4 u5_mult_82_FS_1_U12 ( .A(u5_mult_82_FS_1_n90), .ZN(
        u5_mult_82_FS_1_n11) );
  INV_X4 u5_mult_82_FS_1_U11 ( .A(u5_mult_82_FS_1_n82), .ZN(
        u5_mult_82_FS_1_n10) );
  INV_X4 u5_mult_82_FS_1_U10 ( .A(u5_mult_82_FS_1_n84), .ZN(u5_mult_82_FS_1_n9) );
  INV_X4 u5_mult_82_FS_1_U9 ( .A(u5_mult_82_FS_1_n80), .ZN(u5_mult_82_FS_1_n8)
         );
  INV_X4 u5_mult_82_FS_1_U8 ( .A(u5_mult_82_FS_1_n76), .ZN(u5_mult_82_FS_1_n7)
         );
  INV_X4 u5_mult_82_FS_1_U7 ( .A(u5_mult_82_FS_1_n72), .ZN(u5_mult_82_FS_1_n6)
         );
  INV_X4 u5_mult_82_FS_1_U6 ( .A(u5_mult_82_FS_1_n274), .ZN(u5_mult_82_FS_1_n5) );
  INV_X4 u5_mult_82_FS_1_U5 ( .A(u5_mult_82_FS_1_n272), .ZN(u5_mult_82_FS_1_n4) );
  INV_X4 u5_mult_82_FS_1_U4 ( .A(u5_mult_82_FS_1_n266), .ZN(u5_mult_82_FS_1_n3) );
  AND2_X4 u5_mult_82_FS_1_U3 ( .A1(u5_mult_82_FS_1_n1), .A2(
        u5_mult_82_FS_1_n264), .ZN(u5_N54) );
  OR2_X4 u5_mult_82_FS_1_U2 ( .A1(u5_mult_82_n107), .A2(u5_mult_82_n6), .ZN(
        u5_mult_82_FS_1_n1) );
endmodule

